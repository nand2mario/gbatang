//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9 (64-bit)
//Part Number: GW5AST-LV138PG484AC1/I0
//Device: GW5AST-138B
//Device Version: B
//Created Time: Sun Jun 30 20:30:04 2024

module vram_hi (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb, byte_ena, byte_enb);

output [31:0] douta;
output [31:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [12:0] ada;
input [31:0] dina;
input [12:0] adb;
input [31:0] dinb;
input [3:0] byte_ena;
input [3:0] byte_enb;

wire [15:0] dpb_inst_0_douta;
wire [15:0] dpb_inst_0_doutb;
wire [15:0] dpb_inst_1_douta;
wire [15:0] dpb_inst_1_doutb;
wire [15:0] dpb_inst_2_douta;
wire [15:0] dpb_inst_2_doutb;
wire [15:0] dpb_inst_3_douta;
wire [15:0] dpb_inst_3_doutb;
wire [15:0] dpb_inst_4_douta;
wire [15:0] dpb_inst_4_doutb;
wire [15:0] dpb_inst_5_douta;
wire [15:0] dpb_inst_5_doutb;
wire [15:0] dpb_inst_6_douta;
wire [15:0] dpb_inst_6_doutb;
wire [15:0] dpb_inst_7_douta;
wire [15:0] dpb_inst_7_doutb;
wire [31:16] dpb_inst_8_douta;
wire [31:16] dpb_inst_8_doutb;
wire [31:16] dpb_inst_9_douta;
wire [31:16] dpb_inst_9_doutb;
wire [31:16] dpb_inst_10_douta;
wire [31:16] dpb_inst_10_doutb;
wire [31:16] dpb_inst_11_douta;
wire [31:16] dpb_inst_11_doutb;
wire [31:16] dpb_inst_12_douta;
wire [31:16] dpb_inst_12_doutb;
wire [31:16] dpb_inst_13_douta;
wire [31:16] dpb_inst_13_doutb;
wire [31:16] dpb_inst_14_douta;
wire [31:16] dpb_inst_14_doutb;
wire [31:16] dpb_inst_15_douta;
wire [31:16] dpb_inst_15_doutb;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire dff_q_4;
wire dff_q_5;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_28;
wire mux_o_29;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_42;
wire mux_o_43;
wire mux_o_44;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_60;
wire mux_o_61;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_74;
wire mux_o_75;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_89;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_119;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_123;
wire mux_o_124;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_147;
wire mux_o_148;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_154;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_164;
wire mux_o_165;
wire mux_o_166;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_179;
wire mux_o_180;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_194;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_224;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_245;
wire mux_o_246;
wire mux_o_247;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_252;
wire mux_o_253;
wire mux_o_254;
wire mux_o_255;
wire mux_o_256;
wire mux_o_257;
wire mux_o_259;
wire mux_o_260;
wire mux_o_261;
wire mux_o_262;
wire mux_o_263;
wire mux_o_264;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_269;
wire mux_o_270;
wire mux_o_271;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_276;
wire mux_o_277;
wire mux_o_278;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_284;
wire mux_o_285;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_297;
wire mux_o_298;
wire mux_o_299;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_304;
wire mux_o_305;
wire mux_o_306;
wire mux_o_308;
wire mux_o_309;
wire mux_o_310;
wire mux_o_311;
wire mux_o_312;
wire mux_o_313;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_329;
wire mux_o_330;
wire mux_o_331;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_360;
wire mux_o_361;
wire mux_o_362;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_371;
wire mux_o_372;
wire mux_o_373;
wire mux_o_374;
wire mux_o_375;
wire mux_o_376;
wire mux_o_378;
wire mux_o_379;
wire mux_o_380;
wire mux_o_381;
wire mux_o_382;
wire mux_o_383;
wire mux_o_385;
wire mux_o_386;
wire mux_o_387;
wire mux_o_388;
wire mux_o_389;
wire mux_o_390;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_399;
wire mux_o_400;
wire mux_o_401;
wire mux_o_402;
wire mux_o_403;
wire mux_o_404;
wire mux_o_406;
wire mux_o_407;
wire mux_o_408;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_413;
wire mux_o_414;
wire mux_o_415;
wire mux_o_416;
wire mux_o_417;
wire mux_o_418;
wire mux_o_420;
wire mux_o_421;
wire mux_o_422;
wire mux_o_423;
wire mux_o_424;
wire mux_o_425;
wire mux_o_427;
wire mux_o_428;
wire mux_o_429;
wire mux_o_430;
wire mux_o_431;
wire mux_o_432;
wire mux_o_434;
wire mux_o_435;
wire mux_o_436;
wire mux_o_437;
wire mux_o_438;
wire mux_o_439;
wire mux_o_441;
wire mux_o_442;
wire mux_o_443;
wire mux_o_444;
wire mux_o_445;
wire mux_o_446;
wire cea_w;
wire ceb_w;
wire gw_gnd;

assign cea_w = ~wrea & cea;
assign ceb_w = ~wreb & ceb;
assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA(dpb_inst_0_douta[15:0]),
    .DOB(dpb_inst_0_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_0.READ_MODE0 = 1'b0;
defparam dpb_inst_0.READ_MODE1 = 1'b0;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 16;
defparam dpb_inst_0.BIT_WIDTH_1 = 16;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";

DPB dpb_inst_1 (
    .DOA(dpb_inst_1_douta[15:0]),
    .DOB(dpb_inst_1_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_1.READ_MODE0 = 1'b0;
defparam dpb_inst_1.READ_MODE1 = 1'b0;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 16;
defparam dpb_inst_1.BIT_WIDTH_1 = 16;
defparam dpb_inst_1.BLK_SEL_0 = 3'b001;
defparam dpb_inst_1.BLK_SEL_1 = 3'b001;
defparam dpb_inst_1.RESET_MODE = "SYNC";

DPB dpb_inst_2 (
    .DOA(dpb_inst_2_douta[15:0]),
    .DOB(dpb_inst_2_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_2.READ_MODE0 = 1'b0;
defparam dpb_inst_2.READ_MODE1 = 1'b0;
defparam dpb_inst_2.WRITE_MODE0 = 2'b00;
defparam dpb_inst_2.WRITE_MODE1 = 2'b00;
defparam dpb_inst_2.BIT_WIDTH_0 = 16;
defparam dpb_inst_2.BIT_WIDTH_1 = 16;
defparam dpb_inst_2.BLK_SEL_0 = 3'b010;
defparam dpb_inst_2.BLK_SEL_1 = 3'b010;
defparam dpb_inst_2.RESET_MODE = "SYNC";

DPB dpb_inst_3 (
    .DOA(dpb_inst_3_douta[15:0]),
    .DOB(dpb_inst_3_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_3.READ_MODE0 = 1'b0;
defparam dpb_inst_3.READ_MODE1 = 1'b0;
defparam dpb_inst_3.WRITE_MODE0 = 2'b00;
defparam dpb_inst_3.WRITE_MODE1 = 2'b00;
defparam dpb_inst_3.BIT_WIDTH_0 = 16;
defparam dpb_inst_3.BIT_WIDTH_1 = 16;
defparam dpb_inst_3.BLK_SEL_0 = 3'b011;
defparam dpb_inst_3.BLK_SEL_1 = 3'b011;
defparam dpb_inst_3.RESET_MODE = "SYNC";

DPB dpb_inst_4 (
    .DOA(dpb_inst_4_douta[15:0]),
    .DOB(dpb_inst_4_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_4.READ_MODE0 = 1'b0;
defparam dpb_inst_4.READ_MODE1 = 1'b0;
defparam dpb_inst_4.WRITE_MODE0 = 2'b00;
defparam dpb_inst_4.WRITE_MODE1 = 2'b00;
defparam dpb_inst_4.BIT_WIDTH_0 = 16;
defparam dpb_inst_4.BIT_WIDTH_1 = 16;
defparam dpb_inst_4.BLK_SEL_0 = 3'b100;
defparam dpb_inst_4.BLK_SEL_1 = 3'b100;
defparam dpb_inst_4.RESET_MODE = "SYNC";

DPB dpb_inst_5 (
    .DOA(dpb_inst_5_douta[15:0]),
    .DOB(dpb_inst_5_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_5.READ_MODE0 = 1'b0;
defparam dpb_inst_5.READ_MODE1 = 1'b0;
defparam dpb_inst_5.WRITE_MODE0 = 2'b00;
defparam dpb_inst_5.WRITE_MODE1 = 2'b00;
defparam dpb_inst_5.BIT_WIDTH_0 = 16;
defparam dpb_inst_5.BIT_WIDTH_1 = 16;
defparam dpb_inst_5.BLK_SEL_0 = 3'b101;
defparam dpb_inst_5.BLK_SEL_1 = 3'b101;
defparam dpb_inst_5.RESET_MODE = "SYNC";

DPB dpb_inst_6 (
    .DOA(dpb_inst_6_douta[15:0]),
    .DOB(dpb_inst_6_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_6.READ_MODE0 = 1'b0;
defparam dpb_inst_6.READ_MODE1 = 1'b0;
defparam dpb_inst_6.WRITE_MODE0 = 2'b00;
defparam dpb_inst_6.WRITE_MODE1 = 2'b00;
defparam dpb_inst_6.BIT_WIDTH_0 = 16;
defparam dpb_inst_6.BIT_WIDTH_1 = 16;
defparam dpb_inst_6.BLK_SEL_0 = 3'b110;
defparam dpb_inst_6.BLK_SEL_1 = 3'b110;
defparam dpb_inst_6.RESET_MODE = "SYNC";

DPB dpb_inst_7 (
    .DOA(dpb_inst_7_douta[15:0]),
    .DOB(dpb_inst_7_doutb[15:0]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[1:0]}),
    .DIA(dina[15:0]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[1:0]}),
    .DIB(dinb[15:0])
);

defparam dpb_inst_7.READ_MODE0 = 1'b0;
defparam dpb_inst_7.READ_MODE1 = 1'b0;
defparam dpb_inst_7.WRITE_MODE0 = 2'b00;
defparam dpb_inst_7.WRITE_MODE1 = 2'b00;
defparam dpb_inst_7.BIT_WIDTH_0 = 16;
defparam dpb_inst_7.BIT_WIDTH_1 = 16;
defparam dpb_inst_7.BLK_SEL_0 = 3'b111;
defparam dpb_inst_7.BLK_SEL_1 = 3'b111;
defparam dpb_inst_7.RESET_MODE = "SYNC";

DPB dpb_inst_8 (
    .DOA(dpb_inst_8_douta[31:16]),
    .DOB(dpb_inst_8_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_8.READ_MODE0 = 1'b0;
defparam dpb_inst_8.READ_MODE1 = 1'b0;
defparam dpb_inst_8.WRITE_MODE0 = 2'b00;
defparam dpb_inst_8.WRITE_MODE1 = 2'b00;
defparam dpb_inst_8.BIT_WIDTH_0 = 16;
defparam dpb_inst_8.BIT_WIDTH_1 = 16;
defparam dpb_inst_8.BLK_SEL_0 = 3'b000;
defparam dpb_inst_8.BLK_SEL_1 = 3'b000;
defparam dpb_inst_8.RESET_MODE = "SYNC";

DPB dpb_inst_9 (
    .DOA(dpb_inst_9_douta[31:16]),
    .DOB(dpb_inst_9_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_9.READ_MODE0 = 1'b0;
defparam dpb_inst_9.READ_MODE1 = 1'b0;
defparam dpb_inst_9.WRITE_MODE0 = 2'b00;
defparam dpb_inst_9.WRITE_MODE1 = 2'b00;
defparam dpb_inst_9.BIT_WIDTH_0 = 16;
defparam dpb_inst_9.BIT_WIDTH_1 = 16;
defparam dpb_inst_9.BLK_SEL_0 = 3'b001;
defparam dpb_inst_9.BLK_SEL_1 = 3'b001;
defparam dpb_inst_9.RESET_MODE = "SYNC";

DPB dpb_inst_10 (
    .DOA(dpb_inst_10_douta[31:16]),
    .DOB(dpb_inst_10_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_10.READ_MODE0 = 1'b0;
defparam dpb_inst_10.READ_MODE1 = 1'b0;
defparam dpb_inst_10.WRITE_MODE0 = 2'b00;
defparam dpb_inst_10.WRITE_MODE1 = 2'b00;
defparam dpb_inst_10.BIT_WIDTH_0 = 16;
defparam dpb_inst_10.BIT_WIDTH_1 = 16;
defparam dpb_inst_10.BLK_SEL_0 = 3'b010;
defparam dpb_inst_10.BLK_SEL_1 = 3'b010;
defparam dpb_inst_10.RESET_MODE = "SYNC";

DPB dpb_inst_11 (
    .DOA(dpb_inst_11_douta[31:16]),
    .DOB(dpb_inst_11_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_11.READ_MODE0 = 1'b0;
defparam dpb_inst_11.READ_MODE1 = 1'b0;
defparam dpb_inst_11.WRITE_MODE0 = 2'b00;
defparam dpb_inst_11.WRITE_MODE1 = 2'b00;
defparam dpb_inst_11.BIT_WIDTH_0 = 16;
defparam dpb_inst_11.BIT_WIDTH_1 = 16;
defparam dpb_inst_11.BLK_SEL_0 = 3'b011;
defparam dpb_inst_11.BLK_SEL_1 = 3'b011;
defparam dpb_inst_11.RESET_MODE = "SYNC";

DPB dpb_inst_12 (
    .DOA(dpb_inst_12_douta[31:16]),
    .DOB(dpb_inst_12_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_12.READ_MODE0 = 1'b0;
defparam dpb_inst_12.READ_MODE1 = 1'b0;
defparam dpb_inst_12.WRITE_MODE0 = 2'b00;
defparam dpb_inst_12.WRITE_MODE1 = 2'b00;
defparam dpb_inst_12.BIT_WIDTH_0 = 16;
defparam dpb_inst_12.BIT_WIDTH_1 = 16;
defparam dpb_inst_12.BLK_SEL_0 = 3'b100;
defparam dpb_inst_12.BLK_SEL_1 = 3'b100;
defparam dpb_inst_12.RESET_MODE = "SYNC";

DPB dpb_inst_13 (
    .DOA(dpb_inst_13_douta[31:16]),
    .DOB(dpb_inst_13_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_13.READ_MODE0 = 1'b0;
defparam dpb_inst_13.READ_MODE1 = 1'b0;
defparam dpb_inst_13.WRITE_MODE0 = 2'b00;
defparam dpb_inst_13.WRITE_MODE1 = 2'b00;
defparam dpb_inst_13.BIT_WIDTH_0 = 16;
defparam dpb_inst_13.BIT_WIDTH_1 = 16;
defparam dpb_inst_13.BLK_SEL_0 = 3'b101;
defparam dpb_inst_13.BLK_SEL_1 = 3'b101;
defparam dpb_inst_13.RESET_MODE = "SYNC";

DPB dpb_inst_14 (
    .DOA(dpb_inst_14_douta[31:16]),
    .DOB(dpb_inst_14_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_14.READ_MODE0 = 1'b0;
defparam dpb_inst_14.READ_MODE1 = 1'b0;
defparam dpb_inst_14.WRITE_MODE0 = 2'b00;
defparam dpb_inst_14.WRITE_MODE1 = 2'b00;
defparam dpb_inst_14.BIT_WIDTH_0 = 16;
defparam dpb_inst_14.BIT_WIDTH_1 = 16;
defparam dpb_inst_14.BLK_SEL_0 = 3'b110;
defparam dpb_inst_14.BLK_SEL_1 = 3'b110;
defparam dpb_inst_14.RESET_MODE = "SYNC";

DPB dpb_inst_15 (
    .DOA(dpb_inst_15_douta[31:16]),
    .DOB(dpb_inst_15_doutb[31:16]),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[12],ada[11],ada[10]}),
    .BLKSELB({adb[12],adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,byte_ena[3:2]}),
    .DIA(dina[31:16]),
    .ADB({adb[9:0],gw_gnd,gw_gnd,byte_enb[3:2]}),
    .DIB(dinb[31:16])
);

defparam dpb_inst_15.READ_MODE0 = 1'b0;
defparam dpb_inst_15.READ_MODE1 = 1'b0;
defparam dpb_inst_15.WRITE_MODE0 = 2'b00;
defparam dpb_inst_15.WRITE_MODE1 = 2'b00;
defparam dpb_inst_15.BIT_WIDTH_0 = 16;
defparam dpb_inst_15.BIT_WIDTH_1 = 16;
defparam dpb_inst_15.BLK_SEL_0 = 3'b111;
defparam dpb_inst_15.BLK_SEL_1 = 3'b111;
defparam dpb_inst_15.RESET_MODE = "SYNC";

DFFRE dff_inst_0 (
  .Q(dff_q_0),
  .D(ada[12]),
  .CLK(clka),
  .CE(cea_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_1 (
  .Q(dff_q_1),
  .D(ada[11]),
  .CLK(clka),
  .CE(cea_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_2 (
  .Q(dff_q_2),
  .D(ada[10]),
  .CLK(clka),
  .CE(cea_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_3 (
  .Q(dff_q_3),
  .D(adb[12]),
  .CLK(clkb),
  .CE(ceb_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_4 (
  .Q(dff_q_4),
  .D(adb[11]),
  .CLK(clkb),
  .CE(ceb_w),
  .RESET(gw_gnd)
);
DFFRE dff_inst_5 (
  .Q(dff_q_5),
  .D(adb[10]),
  .CLK(clkb),
  .CE(ceb_w),
  .RESET(gw_gnd)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(dpb_inst_0_douta[0]),
  .I1(dpb_inst_1_douta[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(dpb_inst_2_douta[0]),
  .I1(dpb_inst_3_douta[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(dpb_inst_4_douta[0]),
  .I1(dpb_inst_5_douta[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(dpb_inst_6_douta[0]),
  .I1(dpb_inst_7_douta[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_1)
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(dff_q_1)
);
MUX2 mux_inst_6 (
  .O(douta[0]),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(dff_q_0)
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(dpb_inst_0_douta[1]),
  .I1(dpb_inst_1_douta[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(dpb_inst_2_douta[1]),
  .I1(dpb_inst_3_douta[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(dpb_inst_4_douta[1]),
  .I1(dpb_inst_5_douta[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(dpb_inst_6_douta[1]),
  .I1(dpb_inst_7_douta[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(mux_o_7),
  .I1(mux_o_8),
  .S0(dff_q_1)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(mux_o_9),
  .I1(mux_o_10),
  .S0(dff_q_1)
);
MUX2 mux_inst_13 (
  .O(douta[1]),
  .I0(mux_o_11),
  .I1(mux_o_12),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(dpb_inst_0_douta[2]),
  .I1(dpb_inst_1_douta[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(dpb_inst_2_douta[2]),
  .I1(dpb_inst_3_douta[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(dpb_inst_4_douta[2]),
  .I1(dpb_inst_5_douta[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(dpb_inst_6_douta[2]),
  .I1(dpb_inst_7_douta[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(dff_q_1)
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(dff_q_1)
);
MUX2 mux_inst_20 (
  .O(douta[2]),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(dff_q_0)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(dpb_inst_0_douta[3]),
  .I1(dpb_inst_1_douta[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(dpb_inst_2_douta[3]),
  .I1(dpb_inst_3_douta[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(dpb_inst_4_douta[3]),
  .I1(dpb_inst_5_douta[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(dpb_inst_6_douta[3]),
  .I1(dpb_inst_7_douta[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(mux_o_21),
  .I1(mux_o_22),
  .S0(dff_q_1)
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(mux_o_23),
  .I1(mux_o_24),
  .S0(dff_q_1)
);
MUX2 mux_inst_27 (
  .O(douta[3]),
  .I0(mux_o_25),
  .I1(mux_o_26),
  .S0(dff_q_0)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(dpb_inst_0_douta[4]),
  .I1(dpb_inst_1_douta[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(dpb_inst_2_douta[4]),
  .I1(dpb_inst_3_douta[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(dpb_inst_4_douta[4]),
  .I1(dpb_inst_5_douta[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(dpb_inst_6_douta[4]),
  .I1(dpb_inst_7_douta[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(mux_o_28),
  .I1(mux_o_29),
  .S0(dff_q_1)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(mux_o_30),
  .I1(mux_o_31),
  .S0(dff_q_1)
);
MUX2 mux_inst_34 (
  .O(douta[4]),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(dff_q_0)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(dpb_inst_0_douta[5]),
  .I1(dpb_inst_1_douta[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(dpb_inst_2_douta[5]),
  .I1(dpb_inst_3_douta[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(dpb_inst_4_douta[5]),
  .I1(dpb_inst_5_douta[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(dpb_inst_6_douta[5]),
  .I1(dpb_inst_7_douta[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_35),
  .I1(mux_o_36),
  .S0(dff_q_1)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_37),
  .I1(mux_o_38),
  .S0(dff_q_1)
);
MUX2 mux_inst_41 (
  .O(douta[5]),
  .I0(mux_o_39),
  .I1(mux_o_40),
  .S0(dff_q_0)
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(dpb_inst_0_douta[6]),
  .I1(dpb_inst_1_douta[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(dpb_inst_2_douta[6]),
  .I1(dpb_inst_3_douta[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(dpb_inst_4_douta[6]),
  .I1(dpb_inst_5_douta[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(dpb_inst_6_douta[6]),
  .I1(dpb_inst_7_douta[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(dff_q_1)
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(mux_o_44),
  .I1(mux_o_45),
  .S0(dff_q_1)
);
MUX2 mux_inst_48 (
  .O(douta[6]),
  .I0(mux_o_46),
  .I1(mux_o_47),
  .S0(dff_q_0)
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(dpb_inst_0_douta[7]),
  .I1(dpb_inst_1_douta[7]),
  .S0(dff_q_2)
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(dpb_inst_2_douta[7]),
  .I1(dpb_inst_3_douta[7]),
  .S0(dff_q_2)
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(dpb_inst_4_douta[7]),
  .I1(dpb_inst_5_douta[7]),
  .S0(dff_q_2)
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(dpb_inst_6_douta[7]),
  .I1(dpb_inst_7_douta[7]),
  .S0(dff_q_2)
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(dff_q_1)
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_51),
  .I1(mux_o_52),
  .S0(dff_q_1)
);
MUX2 mux_inst_55 (
  .O(douta[7]),
  .I0(mux_o_53),
  .I1(mux_o_54),
  .S0(dff_q_0)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(dpb_inst_0_douta[8]),
  .I1(dpb_inst_1_douta[8]),
  .S0(dff_q_2)
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(dpb_inst_2_douta[8]),
  .I1(dpb_inst_3_douta[8]),
  .S0(dff_q_2)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(dpb_inst_4_douta[8]),
  .I1(dpb_inst_5_douta[8]),
  .S0(dff_q_2)
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(dpb_inst_6_douta[8]),
  .I1(dpb_inst_7_douta[8]),
  .S0(dff_q_2)
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(mux_o_56),
  .I1(mux_o_57),
  .S0(dff_q_1)
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(mux_o_58),
  .I1(mux_o_59),
  .S0(dff_q_1)
);
MUX2 mux_inst_62 (
  .O(douta[8]),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(dff_q_0)
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(dpb_inst_0_douta[9]),
  .I1(dpb_inst_1_douta[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(dpb_inst_2_douta[9]),
  .I1(dpb_inst_3_douta[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(dpb_inst_4_douta[9]),
  .I1(dpb_inst_5_douta[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(dpb_inst_6_douta[9]),
  .I1(dpb_inst_7_douta[9]),
  .S0(dff_q_2)
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(mux_o_63),
  .I1(mux_o_64),
  .S0(dff_q_1)
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(mux_o_65),
  .I1(mux_o_66),
  .S0(dff_q_1)
);
MUX2 mux_inst_69 (
  .O(douta[9]),
  .I0(mux_o_67),
  .I1(mux_o_68),
  .S0(dff_q_0)
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(dpb_inst_0_douta[10]),
  .I1(dpb_inst_1_douta[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(dpb_inst_2_douta[10]),
  .I1(dpb_inst_3_douta[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(dpb_inst_4_douta[10]),
  .I1(dpb_inst_5_douta[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(dpb_inst_6_douta[10]),
  .I1(dpb_inst_7_douta[10]),
  .S0(dff_q_2)
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(dff_q_1)
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(dff_q_1)
);
MUX2 mux_inst_76 (
  .O(douta[10]),
  .I0(mux_o_74),
  .I1(mux_o_75),
  .S0(dff_q_0)
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(dpb_inst_0_douta[11]),
  .I1(dpb_inst_1_douta[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(dpb_inst_2_douta[11]),
  .I1(dpb_inst_3_douta[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(dpb_inst_4_douta[11]),
  .I1(dpb_inst_5_douta[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(dpb_inst_6_douta[11]),
  .I1(dpb_inst_7_douta[11]),
  .S0(dff_q_2)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(dff_q_1)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(dff_q_1)
);
MUX2 mux_inst_83 (
  .O(douta[11]),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(dff_q_0)
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(dpb_inst_0_douta[12]),
  .I1(dpb_inst_1_douta[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(dpb_inst_2_douta[12]),
  .I1(dpb_inst_3_douta[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(dpb_inst_4_douta[12]),
  .I1(dpb_inst_5_douta[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(dpb_inst_6_douta[12]),
  .I1(dpb_inst_7_douta[12]),
  .S0(dff_q_2)
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(mux_o_84),
  .I1(mux_o_85),
  .S0(dff_q_1)
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(mux_o_86),
  .I1(mux_o_87),
  .S0(dff_q_1)
);
MUX2 mux_inst_90 (
  .O(douta[12]),
  .I0(mux_o_88),
  .I1(mux_o_89),
  .S0(dff_q_0)
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(dpb_inst_0_douta[13]),
  .I1(dpb_inst_1_douta[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(dpb_inst_2_douta[13]),
  .I1(dpb_inst_3_douta[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(dpb_inst_4_douta[13]),
  .I1(dpb_inst_5_douta[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(dpb_inst_6_douta[13]),
  .I1(dpb_inst_7_douta[13]),
  .S0(dff_q_2)
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(mux_o_91),
  .I1(mux_o_92),
  .S0(dff_q_1)
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(mux_o_93),
  .I1(mux_o_94),
  .S0(dff_q_1)
);
MUX2 mux_inst_97 (
  .O(douta[13]),
  .I0(mux_o_95),
  .I1(mux_o_96),
  .S0(dff_q_0)
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(dpb_inst_0_douta[14]),
  .I1(dpb_inst_1_douta[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(dpb_inst_2_douta[14]),
  .I1(dpb_inst_3_douta[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(dpb_inst_4_douta[14]),
  .I1(dpb_inst_5_douta[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(dpb_inst_6_douta[14]),
  .I1(dpb_inst_7_douta[14]),
  .S0(dff_q_2)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_98),
  .I1(mux_o_99),
  .S0(dff_q_1)
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(mux_o_100),
  .I1(mux_o_101),
  .S0(dff_q_1)
);
MUX2 mux_inst_104 (
  .O(douta[14]),
  .I0(mux_o_102),
  .I1(mux_o_103),
  .S0(dff_q_0)
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(dpb_inst_0_douta[15]),
  .I1(dpb_inst_1_douta[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(dpb_inst_2_douta[15]),
  .I1(dpb_inst_3_douta[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(dpb_inst_4_douta[15]),
  .I1(dpb_inst_5_douta[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(dpb_inst_6_douta[15]),
  .I1(dpb_inst_7_douta[15]),
  .S0(dff_q_2)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(mux_o_105),
  .I1(mux_o_106),
  .S0(dff_q_1)
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(dff_q_1)
);
MUX2 mux_inst_111 (
  .O(douta[15]),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(dff_q_0)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(dpb_inst_8_douta[16]),
  .I1(dpb_inst_9_douta[16]),
  .S0(dff_q_2)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(dpb_inst_10_douta[16]),
  .I1(dpb_inst_11_douta[16]),
  .S0(dff_q_2)
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(dpb_inst_12_douta[16]),
  .I1(dpb_inst_13_douta[16]),
  .S0(dff_q_2)
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(dpb_inst_14_douta[16]),
  .I1(dpb_inst_15_douta[16]),
  .S0(dff_q_2)
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_112),
  .I1(mux_o_113),
  .S0(dff_q_1)
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_114),
  .I1(mux_o_115),
  .S0(dff_q_1)
);
MUX2 mux_inst_118 (
  .O(douta[16]),
  .I0(mux_o_116),
  .I1(mux_o_117),
  .S0(dff_q_0)
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(dpb_inst_8_douta[17]),
  .I1(dpb_inst_9_douta[17]),
  .S0(dff_q_2)
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(dpb_inst_10_douta[17]),
  .I1(dpb_inst_11_douta[17]),
  .S0(dff_q_2)
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(dpb_inst_12_douta[17]),
  .I1(dpb_inst_13_douta[17]),
  .S0(dff_q_2)
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(dpb_inst_14_douta[17]),
  .I1(dpb_inst_15_douta[17]),
  .S0(dff_q_2)
);
MUX2 mux_inst_123 (
  .O(mux_o_123),
  .I0(mux_o_119),
  .I1(mux_o_120),
  .S0(dff_q_1)
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(mux_o_121),
  .I1(mux_o_122),
  .S0(dff_q_1)
);
MUX2 mux_inst_125 (
  .O(douta[17]),
  .I0(mux_o_123),
  .I1(mux_o_124),
  .S0(dff_q_0)
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(dpb_inst_8_douta[18]),
  .I1(dpb_inst_9_douta[18]),
  .S0(dff_q_2)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(dpb_inst_10_douta[18]),
  .I1(dpb_inst_11_douta[18]),
  .S0(dff_q_2)
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(dpb_inst_12_douta[18]),
  .I1(dpb_inst_13_douta[18]),
  .S0(dff_q_2)
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(dpb_inst_14_douta[18]),
  .I1(dpb_inst_15_douta[18]),
  .S0(dff_q_2)
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(dff_q_1)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(mux_o_128),
  .I1(mux_o_129),
  .S0(dff_q_1)
);
MUX2 mux_inst_132 (
  .O(douta[18]),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(dff_q_0)
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(dpb_inst_8_douta[19]),
  .I1(dpb_inst_9_douta[19]),
  .S0(dff_q_2)
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(dpb_inst_10_douta[19]),
  .I1(dpb_inst_11_douta[19]),
  .S0(dff_q_2)
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(dpb_inst_12_douta[19]),
  .I1(dpb_inst_13_douta[19]),
  .S0(dff_q_2)
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(dpb_inst_14_douta[19]),
  .I1(dpb_inst_15_douta[19]),
  .S0(dff_q_2)
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(mux_o_133),
  .I1(mux_o_134),
  .S0(dff_q_1)
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(mux_o_135),
  .I1(mux_o_136),
  .S0(dff_q_1)
);
MUX2 mux_inst_139 (
  .O(douta[19]),
  .I0(mux_o_137),
  .I1(mux_o_138),
  .S0(dff_q_0)
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(dpb_inst_8_douta[20]),
  .I1(dpb_inst_9_douta[20]),
  .S0(dff_q_2)
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(dpb_inst_10_douta[20]),
  .I1(dpb_inst_11_douta[20]),
  .S0(dff_q_2)
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(dpb_inst_12_douta[20]),
  .I1(dpb_inst_13_douta[20]),
  .S0(dff_q_2)
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(dpb_inst_14_douta[20]),
  .I1(dpb_inst_15_douta[20]),
  .S0(dff_q_2)
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(mux_o_140),
  .I1(mux_o_141),
  .S0(dff_q_1)
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(mux_o_142),
  .I1(mux_o_143),
  .S0(dff_q_1)
);
MUX2 mux_inst_146 (
  .O(douta[20]),
  .I0(mux_o_144),
  .I1(mux_o_145),
  .S0(dff_q_0)
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(dpb_inst_8_douta[21]),
  .I1(dpb_inst_9_douta[21]),
  .S0(dff_q_2)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(dpb_inst_10_douta[21]),
  .I1(dpb_inst_11_douta[21]),
  .S0(dff_q_2)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(dpb_inst_12_douta[21]),
  .I1(dpb_inst_13_douta[21]),
  .S0(dff_q_2)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(dpb_inst_14_douta[21]),
  .I1(dpb_inst_15_douta[21]),
  .S0(dff_q_2)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(mux_o_147),
  .I1(mux_o_148),
  .S0(dff_q_1)
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(mux_o_149),
  .I1(mux_o_150),
  .S0(dff_q_1)
);
MUX2 mux_inst_153 (
  .O(douta[21]),
  .I0(mux_o_151),
  .I1(mux_o_152),
  .S0(dff_q_0)
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(dpb_inst_8_douta[22]),
  .I1(dpb_inst_9_douta[22]),
  .S0(dff_q_2)
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(dpb_inst_10_douta[22]),
  .I1(dpb_inst_11_douta[22]),
  .S0(dff_q_2)
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(dpb_inst_12_douta[22]),
  .I1(dpb_inst_13_douta[22]),
  .S0(dff_q_2)
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(dpb_inst_14_douta[22]),
  .I1(dpb_inst_15_douta[22]),
  .S0(dff_q_2)
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(mux_o_154),
  .I1(mux_o_155),
  .S0(dff_q_1)
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(mux_o_156),
  .I1(mux_o_157),
  .S0(dff_q_1)
);
MUX2 mux_inst_160 (
  .O(douta[22]),
  .I0(mux_o_158),
  .I1(mux_o_159),
  .S0(dff_q_0)
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(dpb_inst_8_douta[23]),
  .I1(dpb_inst_9_douta[23]),
  .S0(dff_q_2)
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(dpb_inst_10_douta[23]),
  .I1(dpb_inst_11_douta[23]),
  .S0(dff_q_2)
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(dpb_inst_12_douta[23]),
  .I1(dpb_inst_13_douta[23]),
  .S0(dff_q_2)
);
MUX2 mux_inst_164 (
  .O(mux_o_164),
  .I0(dpb_inst_14_douta[23]),
  .I1(dpb_inst_15_douta[23]),
  .S0(dff_q_2)
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(mux_o_161),
  .I1(mux_o_162),
  .S0(dff_q_1)
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(mux_o_163),
  .I1(mux_o_164),
  .S0(dff_q_1)
);
MUX2 mux_inst_167 (
  .O(douta[23]),
  .I0(mux_o_165),
  .I1(mux_o_166),
  .S0(dff_q_0)
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(dpb_inst_8_douta[24]),
  .I1(dpb_inst_9_douta[24]),
  .S0(dff_q_2)
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(dpb_inst_10_douta[24]),
  .I1(dpb_inst_11_douta[24]),
  .S0(dff_q_2)
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(dpb_inst_12_douta[24]),
  .I1(dpb_inst_13_douta[24]),
  .S0(dff_q_2)
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(dpb_inst_14_douta[24]),
  .I1(dpb_inst_15_douta[24]),
  .S0(dff_q_2)
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(mux_o_168),
  .I1(mux_o_169),
  .S0(dff_q_1)
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(mux_o_170),
  .I1(mux_o_171),
  .S0(dff_q_1)
);
MUX2 mux_inst_174 (
  .O(douta[24]),
  .I0(mux_o_172),
  .I1(mux_o_173),
  .S0(dff_q_0)
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(dpb_inst_8_douta[25]),
  .I1(dpb_inst_9_douta[25]),
  .S0(dff_q_2)
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(dpb_inst_10_douta[25]),
  .I1(dpb_inst_11_douta[25]),
  .S0(dff_q_2)
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(dpb_inst_12_douta[25]),
  .I1(dpb_inst_13_douta[25]),
  .S0(dff_q_2)
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(dpb_inst_14_douta[25]),
  .I1(dpb_inst_15_douta[25]),
  .S0(dff_q_2)
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(mux_o_175),
  .I1(mux_o_176),
  .S0(dff_q_1)
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(mux_o_177),
  .I1(mux_o_178),
  .S0(dff_q_1)
);
MUX2 mux_inst_181 (
  .O(douta[25]),
  .I0(mux_o_179),
  .I1(mux_o_180),
  .S0(dff_q_0)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(dpb_inst_8_douta[26]),
  .I1(dpb_inst_9_douta[26]),
  .S0(dff_q_2)
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(dpb_inst_10_douta[26]),
  .I1(dpb_inst_11_douta[26]),
  .S0(dff_q_2)
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(dpb_inst_12_douta[26]),
  .I1(dpb_inst_13_douta[26]),
  .S0(dff_q_2)
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(dpb_inst_14_douta[26]),
  .I1(dpb_inst_15_douta[26]),
  .S0(dff_q_2)
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(mux_o_182),
  .I1(mux_o_183),
  .S0(dff_q_1)
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(mux_o_184),
  .I1(mux_o_185),
  .S0(dff_q_1)
);
MUX2 mux_inst_188 (
  .O(douta[26]),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(dff_q_0)
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(dpb_inst_8_douta[27]),
  .I1(dpb_inst_9_douta[27]),
  .S0(dff_q_2)
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(dpb_inst_10_douta[27]),
  .I1(dpb_inst_11_douta[27]),
  .S0(dff_q_2)
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(dpb_inst_12_douta[27]),
  .I1(dpb_inst_13_douta[27]),
  .S0(dff_q_2)
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(dpb_inst_14_douta[27]),
  .I1(dpb_inst_15_douta[27]),
  .S0(dff_q_2)
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(mux_o_189),
  .I1(mux_o_190),
  .S0(dff_q_1)
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(mux_o_191),
  .I1(mux_o_192),
  .S0(dff_q_1)
);
MUX2 mux_inst_195 (
  .O(douta[27]),
  .I0(mux_o_193),
  .I1(mux_o_194),
  .S0(dff_q_0)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(dpb_inst_8_douta[28]),
  .I1(dpb_inst_9_douta[28]),
  .S0(dff_q_2)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(dpb_inst_10_douta[28]),
  .I1(dpb_inst_11_douta[28]),
  .S0(dff_q_2)
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(dpb_inst_12_douta[28]),
  .I1(dpb_inst_13_douta[28]),
  .S0(dff_q_2)
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(dpb_inst_14_douta[28]),
  .I1(dpb_inst_15_douta[28]),
  .S0(dff_q_2)
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(mux_o_196),
  .I1(mux_o_197),
  .S0(dff_q_1)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(mux_o_198),
  .I1(mux_o_199),
  .S0(dff_q_1)
);
MUX2 mux_inst_202 (
  .O(douta[28]),
  .I0(mux_o_200),
  .I1(mux_o_201),
  .S0(dff_q_0)
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(dpb_inst_8_douta[29]),
  .I1(dpb_inst_9_douta[29]),
  .S0(dff_q_2)
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(dpb_inst_10_douta[29]),
  .I1(dpb_inst_11_douta[29]),
  .S0(dff_q_2)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(dpb_inst_12_douta[29]),
  .I1(dpb_inst_13_douta[29]),
  .S0(dff_q_2)
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(dpb_inst_14_douta[29]),
  .I1(dpb_inst_15_douta[29]),
  .S0(dff_q_2)
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(mux_o_203),
  .I1(mux_o_204),
  .S0(dff_q_1)
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(dff_q_1)
);
MUX2 mux_inst_209 (
  .O(douta[29]),
  .I0(mux_o_207),
  .I1(mux_o_208),
  .S0(dff_q_0)
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(dpb_inst_8_douta[30]),
  .I1(dpb_inst_9_douta[30]),
  .S0(dff_q_2)
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(dpb_inst_10_douta[30]),
  .I1(dpb_inst_11_douta[30]),
  .S0(dff_q_2)
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(dpb_inst_12_douta[30]),
  .I1(dpb_inst_13_douta[30]),
  .S0(dff_q_2)
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(dpb_inst_14_douta[30]),
  .I1(dpb_inst_15_douta[30]),
  .S0(dff_q_2)
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(mux_o_210),
  .I1(mux_o_211),
  .S0(dff_q_1)
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(mux_o_212),
  .I1(mux_o_213),
  .S0(dff_q_1)
);
MUX2 mux_inst_216 (
  .O(douta[30]),
  .I0(mux_o_214),
  .I1(mux_o_215),
  .S0(dff_q_0)
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(dpb_inst_8_douta[31]),
  .I1(dpb_inst_9_douta[31]),
  .S0(dff_q_2)
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(dpb_inst_10_douta[31]),
  .I1(dpb_inst_11_douta[31]),
  .S0(dff_q_2)
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(dpb_inst_12_douta[31]),
  .I1(dpb_inst_13_douta[31]),
  .S0(dff_q_2)
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(dpb_inst_14_douta[31]),
  .I1(dpb_inst_15_douta[31]),
  .S0(dff_q_2)
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(mux_o_217),
  .I1(mux_o_218),
  .S0(dff_q_1)
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(mux_o_219),
  .I1(mux_o_220),
  .S0(dff_q_1)
);
MUX2 mux_inst_223 (
  .O(douta[31]),
  .I0(mux_o_221),
  .I1(mux_o_222),
  .S0(dff_q_0)
);
MUX2 mux_inst_224 (
  .O(mux_o_224),
  .I0(dpb_inst_0_doutb[0]),
  .I1(dpb_inst_1_doutb[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(dpb_inst_2_doutb[0]),
  .I1(dpb_inst_3_doutb[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(dpb_inst_4_doutb[0]),
  .I1(dpb_inst_5_doutb[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(dpb_inst_6_doutb[0]),
  .I1(dpb_inst_7_doutb[0]),
  .S0(dff_q_5)
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(mux_o_224),
  .I1(mux_o_225),
  .S0(dff_q_4)
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(mux_o_226),
  .I1(mux_o_227),
  .S0(dff_q_4)
);
MUX2 mux_inst_230 (
  .O(doutb[0]),
  .I0(mux_o_228),
  .I1(mux_o_229),
  .S0(dff_q_3)
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(dpb_inst_0_doutb[1]),
  .I1(dpb_inst_1_doutb[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(dpb_inst_2_doutb[1]),
  .I1(dpb_inst_3_doutb[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(dpb_inst_4_doutb[1]),
  .I1(dpb_inst_5_doutb[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(dpb_inst_6_doutb[1]),
  .I1(dpb_inst_7_doutb[1]),
  .S0(dff_q_5)
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(dff_q_4)
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(dff_q_4)
);
MUX2 mux_inst_237 (
  .O(doutb[1]),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(dff_q_3)
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(dpb_inst_0_doutb[2]),
  .I1(dpb_inst_1_doutb[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(dpb_inst_2_doutb[2]),
  .I1(dpb_inst_3_doutb[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(dpb_inst_4_doutb[2]),
  .I1(dpb_inst_5_doutb[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(dpb_inst_6_doutb[2]),
  .I1(dpb_inst_7_doutb[2]),
  .S0(dff_q_5)
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(mux_o_238),
  .I1(mux_o_239),
  .S0(dff_q_4)
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(mux_o_240),
  .I1(mux_o_241),
  .S0(dff_q_4)
);
MUX2 mux_inst_244 (
  .O(doutb[2]),
  .I0(mux_o_242),
  .I1(mux_o_243),
  .S0(dff_q_3)
);
MUX2 mux_inst_245 (
  .O(mux_o_245),
  .I0(dpb_inst_0_doutb[3]),
  .I1(dpb_inst_1_doutb[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(dpb_inst_2_doutb[3]),
  .I1(dpb_inst_3_doutb[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(dpb_inst_4_doutb[3]),
  .I1(dpb_inst_5_doutb[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(dpb_inst_6_doutb[3]),
  .I1(dpb_inst_7_doutb[3]),
  .S0(dff_q_5)
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(mux_o_245),
  .I1(mux_o_246),
  .S0(dff_q_4)
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(mux_o_247),
  .I1(mux_o_248),
  .S0(dff_q_4)
);
MUX2 mux_inst_251 (
  .O(doutb[3]),
  .I0(mux_o_249),
  .I1(mux_o_250),
  .S0(dff_q_3)
);
MUX2 mux_inst_252 (
  .O(mux_o_252),
  .I0(dpb_inst_0_doutb[4]),
  .I1(dpb_inst_1_doutb[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(dpb_inst_2_doutb[4]),
  .I1(dpb_inst_3_doutb[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_254 (
  .O(mux_o_254),
  .I0(dpb_inst_4_doutb[4]),
  .I1(dpb_inst_5_doutb[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(dpb_inst_6_doutb[4]),
  .I1(dpb_inst_7_doutb[4]),
  .S0(dff_q_5)
);
MUX2 mux_inst_256 (
  .O(mux_o_256),
  .I0(mux_o_252),
  .I1(mux_o_253),
  .S0(dff_q_4)
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(mux_o_254),
  .I1(mux_o_255),
  .S0(dff_q_4)
);
MUX2 mux_inst_258 (
  .O(doutb[4]),
  .I0(mux_o_256),
  .I1(mux_o_257),
  .S0(dff_q_3)
);
MUX2 mux_inst_259 (
  .O(mux_o_259),
  .I0(dpb_inst_0_doutb[5]),
  .I1(dpb_inst_1_doutb[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(dpb_inst_2_doutb[5]),
  .I1(dpb_inst_3_doutb[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(dpb_inst_4_doutb[5]),
  .I1(dpb_inst_5_doutb[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_262 (
  .O(mux_o_262),
  .I0(dpb_inst_6_doutb[5]),
  .I1(dpb_inst_7_doutb[5]),
  .S0(dff_q_5)
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(mux_o_259),
  .I1(mux_o_260),
  .S0(dff_q_4)
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(mux_o_261),
  .I1(mux_o_262),
  .S0(dff_q_4)
);
MUX2 mux_inst_265 (
  .O(doutb[5]),
  .I0(mux_o_263),
  .I1(mux_o_264),
  .S0(dff_q_3)
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(dpb_inst_0_doutb[6]),
  .I1(dpb_inst_1_doutb[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(dpb_inst_2_doutb[6]),
  .I1(dpb_inst_3_doutb[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(dpb_inst_4_doutb[6]),
  .I1(dpb_inst_5_doutb[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_269 (
  .O(mux_o_269),
  .I0(dpb_inst_6_doutb[6]),
  .I1(dpb_inst_7_doutb[6]),
  .S0(dff_q_5)
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(mux_o_266),
  .I1(mux_o_267),
  .S0(dff_q_4)
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(mux_o_268),
  .I1(mux_o_269),
  .S0(dff_q_4)
);
MUX2 mux_inst_272 (
  .O(doutb[6]),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(dff_q_3)
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(dpb_inst_0_doutb[7]),
  .I1(dpb_inst_1_doutb[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(dpb_inst_2_doutb[7]),
  .I1(dpb_inst_3_doutb[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(dpb_inst_4_doutb[7]),
  .I1(dpb_inst_5_doutb[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_276 (
  .O(mux_o_276),
  .I0(dpb_inst_6_doutb[7]),
  .I1(dpb_inst_7_doutb[7]),
  .S0(dff_q_5)
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(mux_o_273),
  .I1(mux_o_274),
  .S0(dff_q_4)
);
MUX2 mux_inst_278 (
  .O(mux_o_278),
  .I0(mux_o_275),
  .I1(mux_o_276),
  .S0(dff_q_4)
);
MUX2 mux_inst_279 (
  .O(doutb[7]),
  .I0(mux_o_277),
  .I1(mux_o_278),
  .S0(dff_q_3)
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(dpb_inst_0_doutb[8]),
  .I1(dpb_inst_1_doutb[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(dpb_inst_2_doutb[8]),
  .I1(dpb_inst_3_doutb[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(dpb_inst_4_doutb[8]),
  .I1(dpb_inst_5_doutb[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(dpb_inst_6_doutb[8]),
  .I1(dpb_inst_7_doutb[8]),
  .S0(dff_q_5)
);
MUX2 mux_inst_284 (
  .O(mux_o_284),
  .I0(mux_o_280),
  .I1(mux_o_281),
  .S0(dff_q_4)
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(mux_o_282),
  .I1(mux_o_283),
  .S0(dff_q_4)
);
MUX2 mux_inst_286 (
  .O(doutb[8]),
  .I0(mux_o_284),
  .I1(mux_o_285),
  .S0(dff_q_3)
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(dpb_inst_0_doutb[9]),
  .I1(dpb_inst_1_doutb[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(dpb_inst_2_doutb[9]),
  .I1(dpb_inst_3_doutb[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(dpb_inst_4_doutb[9]),
  .I1(dpb_inst_5_doutb[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(dpb_inst_6_doutb[9]),
  .I1(dpb_inst_7_doutb[9]),
  .S0(dff_q_5)
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(mux_o_287),
  .I1(mux_o_288),
  .S0(dff_q_4)
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(mux_o_289),
  .I1(mux_o_290),
  .S0(dff_q_4)
);
MUX2 mux_inst_293 (
  .O(doutb[9]),
  .I0(mux_o_291),
  .I1(mux_o_292),
  .S0(dff_q_3)
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(dpb_inst_0_doutb[10]),
  .I1(dpb_inst_1_doutb[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(dpb_inst_2_doutb[10]),
  .I1(dpb_inst_3_doutb[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(dpb_inst_4_doutb[10]),
  .I1(dpb_inst_5_doutb[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_297 (
  .O(mux_o_297),
  .I0(dpb_inst_6_doutb[10]),
  .I1(dpb_inst_7_doutb[10]),
  .S0(dff_q_5)
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(mux_o_294),
  .I1(mux_o_295),
  .S0(dff_q_4)
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(mux_o_296),
  .I1(mux_o_297),
  .S0(dff_q_4)
);
MUX2 mux_inst_300 (
  .O(doutb[10]),
  .I0(mux_o_298),
  .I1(mux_o_299),
  .S0(dff_q_3)
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(dpb_inst_0_doutb[11]),
  .I1(dpb_inst_1_doutb[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(dpb_inst_2_doutb[11]),
  .I1(dpb_inst_3_doutb[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(dpb_inst_4_doutb[11]),
  .I1(dpb_inst_5_doutb[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_304 (
  .O(mux_o_304),
  .I0(dpb_inst_6_doutb[11]),
  .I1(dpb_inst_7_doutb[11]),
  .S0(dff_q_5)
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(mux_o_301),
  .I1(mux_o_302),
  .S0(dff_q_4)
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(mux_o_303),
  .I1(mux_o_304),
  .S0(dff_q_4)
);
MUX2 mux_inst_307 (
  .O(doutb[11]),
  .I0(mux_o_305),
  .I1(mux_o_306),
  .S0(dff_q_3)
);
MUX2 mux_inst_308 (
  .O(mux_o_308),
  .I0(dpb_inst_0_doutb[12]),
  .I1(dpb_inst_1_doutb[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(dpb_inst_2_doutb[12]),
  .I1(dpb_inst_3_doutb[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(dpb_inst_4_doutb[12]),
  .I1(dpb_inst_5_doutb[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_311 (
  .O(mux_o_311),
  .I0(dpb_inst_6_doutb[12]),
  .I1(dpb_inst_7_doutb[12]),
  .S0(dff_q_5)
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(mux_o_308),
  .I1(mux_o_309),
  .S0(dff_q_4)
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(mux_o_310),
  .I1(mux_o_311),
  .S0(dff_q_4)
);
MUX2 mux_inst_314 (
  .O(doutb[12]),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(dff_q_3)
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(dpb_inst_0_doutb[13]),
  .I1(dpb_inst_1_doutb[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(dpb_inst_2_doutb[13]),
  .I1(dpb_inst_3_doutb[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(dpb_inst_4_doutb[13]),
  .I1(dpb_inst_5_doutb[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(dpb_inst_6_doutb[13]),
  .I1(dpb_inst_7_doutb[13]),
  .S0(dff_q_5)
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(mux_o_315),
  .I1(mux_o_316),
  .S0(dff_q_4)
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(mux_o_317),
  .I1(mux_o_318),
  .S0(dff_q_4)
);
MUX2 mux_inst_321 (
  .O(doutb[13]),
  .I0(mux_o_319),
  .I1(mux_o_320),
  .S0(dff_q_3)
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(dpb_inst_0_doutb[14]),
  .I1(dpb_inst_1_doutb[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(dpb_inst_2_doutb[14]),
  .I1(dpb_inst_3_doutb[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(dpb_inst_4_doutb[14]),
  .I1(dpb_inst_5_doutb[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(dpb_inst_6_doutb[14]),
  .I1(dpb_inst_7_doutb[14]),
  .S0(dff_q_5)
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(mux_o_322),
  .I1(mux_o_323),
  .S0(dff_q_4)
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(mux_o_324),
  .I1(mux_o_325),
  .S0(dff_q_4)
);
MUX2 mux_inst_328 (
  .O(doutb[14]),
  .I0(mux_o_326),
  .I1(mux_o_327),
  .S0(dff_q_3)
);
MUX2 mux_inst_329 (
  .O(mux_o_329),
  .I0(dpb_inst_0_doutb[15]),
  .I1(dpb_inst_1_doutb[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(dpb_inst_2_doutb[15]),
  .I1(dpb_inst_3_doutb[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(dpb_inst_4_doutb[15]),
  .I1(dpb_inst_5_doutb[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(dpb_inst_6_doutb[15]),
  .I1(dpb_inst_7_doutb[15]),
  .S0(dff_q_5)
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(mux_o_329),
  .I1(mux_o_330),
  .S0(dff_q_4)
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(mux_o_331),
  .I1(mux_o_332),
  .S0(dff_q_4)
);
MUX2 mux_inst_335 (
  .O(doutb[15]),
  .I0(mux_o_333),
  .I1(mux_o_334),
  .S0(dff_q_3)
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(dpb_inst_8_doutb[16]),
  .I1(dpb_inst_9_doutb[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(dpb_inst_10_doutb[16]),
  .I1(dpb_inst_11_doutb[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(dpb_inst_12_doutb[16]),
  .I1(dpb_inst_13_doutb[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(dpb_inst_14_doutb[16]),
  .I1(dpb_inst_15_doutb[16]),
  .S0(dff_q_5)
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(mux_o_336),
  .I1(mux_o_337),
  .S0(dff_q_4)
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(mux_o_338),
  .I1(mux_o_339),
  .S0(dff_q_4)
);
MUX2 mux_inst_342 (
  .O(doutb[16]),
  .I0(mux_o_340),
  .I1(mux_o_341),
  .S0(dff_q_3)
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(dpb_inst_8_doutb[17]),
  .I1(dpb_inst_9_doutb[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(dpb_inst_10_doutb[17]),
  .I1(dpb_inst_11_doutb[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(dpb_inst_12_doutb[17]),
  .I1(dpb_inst_13_doutb[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(dpb_inst_14_doutb[17]),
  .I1(dpb_inst_15_doutb[17]),
  .S0(dff_q_5)
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(mux_o_343),
  .I1(mux_o_344),
  .S0(dff_q_4)
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(mux_o_345),
  .I1(mux_o_346),
  .S0(dff_q_4)
);
MUX2 mux_inst_349 (
  .O(doutb[17]),
  .I0(mux_o_347),
  .I1(mux_o_348),
  .S0(dff_q_3)
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(dpb_inst_8_doutb[18]),
  .I1(dpb_inst_9_doutb[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(dpb_inst_10_doutb[18]),
  .I1(dpb_inst_11_doutb[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(dpb_inst_12_doutb[18]),
  .I1(dpb_inst_13_doutb[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(dpb_inst_14_doutb[18]),
  .I1(dpb_inst_15_doutb[18]),
  .S0(dff_q_5)
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(mux_o_350),
  .I1(mux_o_351),
  .S0(dff_q_4)
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(mux_o_352),
  .I1(mux_o_353),
  .S0(dff_q_4)
);
MUX2 mux_inst_356 (
  .O(doutb[18]),
  .I0(mux_o_354),
  .I1(mux_o_355),
  .S0(dff_q_3)
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(dpb_inst_8_doutb[19]),
  .I1(dpb_inst_9_doutb[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(dpb_inst_10_doutb[19]),
  .I1(dpb_inst_11_doutb[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(dpb_inst_12_doutb[19]),
  .I1(dpb_inst_13_doutb[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_360 (
  .O(mux_o_360),
  .I0(dpb_inst_14_doutb[19]),
  .I1(dpb_inst_15_doutb[19]),
  .S0(dff_q_5)
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(mux_o_357),
  .I1(mux_o_358),
  .S0(dff_q_4)
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(mux_o_359),
  .I1(mux_o_360),
  .S0(dff_q_4)
);
MUX2 mux_inst_363 (
  .O(doutb[19]),
  .I0(mux_o_361),
  .I1(mux_o_362),
  .S0(dff_q_3)
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(dpb_inst_8_doutb[20]),
  .I1(dpb_inst_9_doutb[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(dpb_inst_10_doutb[20]),
  .I1(dpb_inst_11_doutb[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(dpb_inst_12_doutb[20]),
  .I1(dpb_inst_13_doutb[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(dpb_inst_14_doutb[20]),
  .I1(dpb_inst_15_doutb[20]),
  .S0(dff_q_5)
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(mux_o_364),
  .I1(mux_o_365),
  .S0(dff_q_4)
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(mux_o_366),
  .I1(mux_o_367),
  .S0(dff_q_4)
);
MUX2 mux_inst_370 (
  .O(doutb[20]),
  .I0(mux_o_368),
  .I1(mux_o_369),
  .S0(dff_q_3)
);
MUX2 mux_inst_371 (
  .O(mux_o_371),
  .I0(dpb_inst_8_doutb[21]),
  .I1(dpb_inst_9_doutb[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(dpb_inst_10_doutb[21]),
  .I1(dpb_inst_11_doutb[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(dpb_inst_12_doutb[21]),
  .I1(dpb_inst_13_doutb[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_374 (
  .O(mux_o_374),
  .I0(dpb_inst_14_doutb[21]),
  .I1(dpb_inst_15_doutb[21]),
  .S0(dff_q_5)
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(mux_o_371),
  .I1(mux_o_372),
  .S0(dff_q_4)
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(mux_o_373),
  .I1(mux_o_374),
  .S0(dff_q_4)
);
MUX2 mux_inst_377 (
  .O(doutb[21]),
  .I0(mux_o_375),
  .I1(mux_o_376),
  .S0(dff_q_3)
);
MUX2 mux_inst_378 (
  .O(mux_o_378),
  .I0(dpb_inst_8_doutb[22]),
  .I1(dpb_inst_9_doutb[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_379 (
  .O(mux_o_379),
  .I0(dpb_inst_10_doutb[22]),
  .I1(dpb_inst_11_doutb[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_380 (
  .O(mux_o_380),
  .I0(dpb_inst_12_doutb[22]),
  .I1(dpb_inst_13_doutb[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_381 (
  .O(mux_o_381),
  .I0(dpb_inst_14_doutb[22]),
  .I1(dpb_inst_15_doutb[22]),
  .S0(dff_q_5)
);
MUX2 mux_inst_382 (
  .O(mux_o_382),
  .I0(mux_o_378),
  .I1(mux_o_379),
  .S0(dff_q_4)
);
MUX2 mux_inst_383 (
  .O(mux_o_383),
  .I0(mux_o_380),
  .I1(mux_o_381),
  .S0(dff_q_4)
);
MUX2 mux_inst_384 (
  .O(doutb[22]),
  .I0(mux_o_382),
  .I1(mux_o_383),
  .S0(dff_q_3)
);
MUX2 mux_inst_385 (
  .O(mux_o_385),
  .I0(dpb_inst_8_doutb[23]),
  .I1(dpb_inst_9_doutb[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_386 (
  .O(mux_o_386),
  .I0(dpb_inst_10_doutb[23]),
  .I1(dpb_inst_11_doutb[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_387 (
  .O(mux_o_387),
  .I0(dpb_inst_12_doutb[23]),
  .I1(dpb_inst_13_doutb[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_388 (
  .O(mux_o_388),
  .I0(dpb_inst_14_doutb[23]),
  .I1(dpb_inst_15_doutb[23]),
  .S0(dff_q_5)
);
MUX2 mux_inst_389 (
  .O(mux_o_389),
  .I0(mux_o_385),
  .I1(mux_o_386),
  .S0(dff_q_4)
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(mux_o_387),
  .I1(mux_o_388),
  .S0(dff_q_4)
);
MUX2 mux_inst_391 (
  .O(doutb[23]),
  .I0(mux_o_389),
  .I1(mux_o_390),
  .S0(dff_q_3)
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(dpb_inst_8_doutb[24]),
  .I1(dpb_inst_9_doutb[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(dpb_inst_10_doutb[24]),
  .I1(dpb_inst_11_doutb[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(dpb_inst_12_doutb[24]),
  .I1(dpb_inst_13_doutb[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(dpb_inst_14_doutb[24]),
  .I1(dpb_inst_15_doutb[24]),
  .S0(dff_q_5)
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(mux_o_392),
  .I1(mux_o_393),
  .S0(dff_q_4)
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(mux_o_394),
  .I1(mux_o_395),
  .S0(dff_q_4)
);
MUX2 mux_inst_398 (
  .O(doutb[24]),
  .I0(mux_o_396),
  .I1(mux_o_397),
  .S0(dff_q_3)
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(dpb_inst_8_doutb[25]),
  .I1(dpb_inst_9_doutb[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(dpb_inst_10_doutb[25]),
  .I1(dpb_inst_11_doutb[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_401 (
  .O(mux_o_401),
  .I0(dpb_inst_12_doutb[25]),
  .I1(dpb_inst_13_doutb[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_402 (
  .O(mux_o_402),
  .I0(dpb_inst_14_doutb[25]),
  .I1(dpb_inst_15_doutb[25]),
  .S0(dff_q_5)
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(mux_o_399),
  .I1(mux_o_400),
  .S0(dff_q_4)
);
MUX2 mux_inst_404 (
  .O(mux_o_404),
  .I0(mux_o_401),
  .I1(mux_o_402),
  .S0(dff_q_4)
);
MUX2 mux_inst_405 (
  .O(doutb[25]),
  .I0(mux_o_403),
  .I1(mux_o_404),
  .S0(dff_q_3)
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(dpb_inst_8_doutb[26]),
  .I1(dpb_inst_9_doutb[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(dpb_inst_10_doutb[26]),
  .I1(dpb_inst_11_doutb[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_408 (
  .O(mux_o_408),
  .I0(dpb_inst_12_doutb[26]),
  .I1(dpb_inst_13_doutb[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(dpb_inst_14_doutb[26]),
  .I1(dpb_inst_15_doutb[26]),
  .S0(dff_q_5)
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(mux_o_406),
  .I1(mux_o_407),
  .S0(dff_q_4)
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(mux_o_408),
  .I1(mux_o_409),
  .S0(dff_q_4)
);
MUX2 mux_inst_412 (
  .O(doutb[26]),
  .I0(mux_o_410),
  .I1(mux_o_411),
  .S0(dff_q_3)
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(dpb_inst_8_doutb[27]),
  .I1(dpb_inst_9_doutb[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(dpb_inst_10_doutb[27]),
  .I1(dpb_inst_11_doutb[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_415 (
  .O(mux_o_415),
  .I0(dpb_inst_12_doutb[27]),
  .I1(dpb_inst_13_doutb[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_416 (
  .O(mux_o_416),
  .I0(dpb_inst_14_doutb[27]),
  .I1(dpb_inst_15_doutb[27]),
  .S0(dff_q_5)
);
MUX2 mux_inst_417 (
  .O(mux_o_417),
  .I0(mux_o_413),
  .I1(mux_o_414),
  .S0(dff_q_4)
);
MUX2 mux_inst_418 (
  .O(mux_o_418),
  .I0(mux_o_415),
  .I1(mux_o_416),
  .S0(dff_q_4)
);
MUX2 mux_inst_419 (
  .O(doutb[27]),
  .I0(mux_o_417),
  .I1(mux_o_418),
  .S0(dff_q_3)
);
MUX2 mux_inst_420 (
  .O(mux_o_420),
  .I0(dpb_inst_8_doutb[28]),
  .I1(dpb_inst_9_doutb[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_421 (
  .O(mux_o_421),
  .I0(dpb_inst_10_doutb[28]),
  .I1(dpb_inst_11_doutb[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_422 (
  .O(mux_o_422),
  .I0(dpb_inst_12_doutb[28]),
  .I1(dpb_inst_13_doutb[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_423 (
  .O(mux_o_423),
  .I0(dpb_inst_14_doutb[28]),
  .I1(dpb_inst_15_doutb[28]),
  .S0(dff_q_5)
);
MUX2 mux_inst_424 (
  .O(mux_o_424),
  .I0(mux_o_420),
  .I1(mux_o_421),
  .S0(dff_q_4)
);
MUX2 mux_inst_425 (
  .O(mux_o_425),
  .I0(mux_o_422),
  .I1(mux_o_423),
  .S0(dff_q_4)
);
MUX2 mux_inst_426 (
  .O(doutb[28]),
  .I0(mux_o_424),
  .I1(mux_o_425),
  .S0(dff_q_3)
);
MUX2 mux_inst_427 (
  .O(mux_o_427),
  .I0(dpb_inst_8_doutb[29]),
  .I1(dpb_inst_9_doutb[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_428 (
  .O(mux_o_428),
  .I0(dpb_inst_10_doutb[29]),
  .I1(dpb_inst_11_doutb[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_429 (
  .O(mux_o_429),
  .I0(dpb_inst_12_doutb[29]),
  .I1(dpb_inst_13_doutb[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_430 (
  .O(mux_o_430),
  .I0(dpb_inst_14_doutb[29]),
  .I1(dpb_inst_15_doutb[29]),
  .S0(dff_q_5)
);
MUX2 mux_inst_431 (
  .O(mux_o_431),
  .I0(mux_o_427),
  .I1(mux_o_428),
  .S0(dff_q_4)
);
MUX2 mux_inst_432 (
  .O(mux_o_432),
  .I0(mux_o_429),
  .I1(mux_o_430),
  .S0(dff_q_4)
);
MUX2 mux_inst_433 (
  .O(doutb[29]),
  .I0(mux_o_431),
  .I1(mux_o_432),
  .S0(dff_q_3)
);
MUX2 mux_inst_434 (
  .O(mux_o_434),
  .I0(dpb_inst_8_doutb[30]),
  .I1(dpb_inst_9_doutb[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_435 (
  .O(mux_o_435),
  .I0(dpb_inst_10_doutb[30]),
  .I1(dpb_inst_11_doutb[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_436 (
  .O(mux_o_436),
  .I0(dpb_inst_12_doutb[30]),
  .I1(dpb_inst_13_doutb[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_437 (
  .O(mux_o_437),
  .I0(dpb_inst_14_doutb[30]),
  .I1(dpb_inst_15_doutb[30]),
  .S0(dff_q_5)
);
MUX2 mux_inst_438 (
  .O(mux_o_438),
  .I0(mux_o_434),
  .I1(mux_o_435),
  .S0(dff_q_4)
);
MUX2 mux_inst_439 (
  .O(mux_o_439),
  .I0(mux_o_436),
  .I1(mux_o_437),
  .S0(dff_q_4)
);
MUX2 mux_inst_440 (
  .O(doutb[30]),
  .I0(mux_o_438),
  .I1(mux_o_439),
  .S0(dff_q_3)
);
MUX2 mux_inst_441 (
  .O(mux_o_441),
  .I0(dpb_inst_8_doutb[31]),
  .I1(dpb_inst_9_doutb[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_442 (
  .O(mux_o_442),
  .I0(dpb_inst_10_doutb[31]),
  .I1(dpb_inst_11_doutb[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_443 (
  .O(mux_o_443),
  .I0(dpb_inst_12_doutb[31]),
  .I1(dpb_inst_13_doutb[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_444 (
  .O(mux_o_444),
  .I0(dpb_inst_14_doutb[31]),
  .I1(dpb_inst_15_doutb[31]),
  .S0(dff_q_5)
);
MUX2 mux_inst_445 (
  .O(mux_o_445),
  .I0(mux_o_441),
  .I1(mux_o_442),
  .S0(dff_q_4)
);
MUX2 mux_inst_446 (
  .O(mux_o_446),
  .I0(mux_o_443),
  .I1(mux_o_444),
  .S0(dff_q_4)
);
MUX2 mux_inst_447 (
  .O(doutb[31]),
  .I0(mux_o_445),
  .I1(mux_o_446),
  .S0(dff_q_3)
);
endmodule //vram_hi

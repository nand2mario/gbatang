`ifndef gba_bios
`define gba_bios

// open source GBA BIOS

// define this to skip logo drawing and go directly to ROM start
`define NO_LOGO

localparam [31:0] GBA_BIOS [0:4095] = '{
    32'hEA00000C,
    32'hEA000015,
    32'hEA000015,
    32'hEA000013,
    32'hEA000012,
    32'hEA000011,
    32'hEA000000,
    32'hEAFFFFFF,
    32'hE92D500F,
    32'hE3A00301,
    32'hE1A0E00F,
    32'hE510F004,
    32'hE8BD500F,
    32'hE25EF004,
    32'hE3A000DF,
    32'hE129F000,
    32'hE3A03301,
    32'hE5C33208,
    32'hEB0005F8,
    32'hE3A02001,
    32'hE5C32208,
    32'hE59F0104,   // 54: ldr	r0, [pc, #260]	        @ 0x160 =DrawLogo
    32'hE59FE104,   // 58: ldr	lr, [pc, #260]	        @ 0x164 =swi_SoftReset
    32'hE12FFF10,   // 5C: bx	r0                      @ draw logo, then link to soft reset
    32'hEAFFFFFE,
    32'hE92D5800,
    32'hE55EC002,
    32'hE28FB03C,
    32'hE79BC10C,
    32'hE14FB000,
    32'hE92D0800,
    32'hE20BB080,
    32'hE38BB01F,
    32'hE129F00B,
    32'hE92D400C,
    32'hE28FE000,
    32'hE12FFF1C,
    32'hE8BD400C,
    32'hE3A0C0D3,
    32'hE129F00C,
    32'hE8BD0800,
    32'hE169F00B,
    32'hE8BD5800,
    32'hE1B0F00E,
    32'h00001804,
    32'h00001524,
    32'h000003D8,
    32'h000003E8,
    32'h00000434,
    32'h000004D4,
    32'h000017A8,
    32'h00001798,
    32'h000004E0,
    32'h000004E4,
    32'h0000056C,
    32'h00000614,
    32'h00000720,
    32'h000007D8,
    32'h000007E4,
    32'h000008E0,
    32'h00000984,
    32'h00000A44,
    32'h00000CDC,
    32'h00000CE4,
    32'h00000F18,
    32'h00000FBC,
    32'h000010C0,
    32'h0000111C,
    32'h000011AC,
    32'h0000015C,
    32'h0000015C,
    32'h0000015C,
    32'h0000015C,
    32'h0000015C,
    32'h0000015C,
    32'h00001218,
    32'h0000015C,
    32'h0000015C,
    32'h0000015C,
    32'h00001500,
    32'h00001504,
    32'h0000015C,
    32'h0000015C,
    32'h000003CC,
    32'h0000015C,
    32'h0000015C,
    32'h00001508,
    32'hE12FFF1E,
`ifdef NO_LOGO
    32'h08000000,   // 160: skip DrawLogo and go directly to ROM start
    // 32'h00001804,   // 160: replace DrawLogo with SoftReset, which goes to ROM start
`else
    32'h000001B8,   // 160: =DrawLogo
`endif
    32'h00001804,   // 164: =swi_SoftReset
    32'hE1A00000,
    32'hE1A00000,
    32'hE0832190,
    32'hE1A00003,
    32'hE12FFF1E,
    32'hE3520000,
    32'h012FFF1E,
    32'hE1A03000,
    32'hE0631001,
    32'hE0800082,
    32'hE3E0C4F1,
    32'hE153000C,
    32'h91D320B0,
    32'h859F2010,
    32'hE18120B3,
    32'hE2833002,
    32'hE1530000,
    32'h1AFFFFF8,
    32'hE12FFF1E,
    32'h00001CAD,
    32'hE92D4008,
    32'hE59FE09C,
    32'hE59FC09C,
    32'hE1A0200E,
    32'hE3A03405,
    32'hE3E004F1,
    32'hE1520000,
    32'h908E1003,
    32'h928114FB,
    32'h91D110B0,
    32'h859F1080,
    32'hE0C310B2,
    32'hE153000C,
    32'hE2822002,
    32'h1AFFFFF6,
    32'hE59F0070,
    32'hE3A01406,
    32'hE3A02000,
    32'hEB000255,
    32'hE59F1064,
    32'hE3A02000,
    32'hE59F0060,
    32'hEB000251,
    32'hE3A03301,
    32'hE3A02C1E,
    32'hE1C320B8,
    32'hE3A02C01,
    32'hE5832000,
    32'hE3A01077,
    32'hE1D320B6,
    32'hE352009F,
    32'h8AFFFFFC,
    32'hE1D320B6,
    32'hE352009F,
    32'h9AFFFFFC,
    32'hE3510000,
    32'hE2411001,
    32'h1AFFFFF6,
    32'hE3A000FF,
    32'hEB0004B2,
    32'hE8BD4008,
    32'hE12FFF1E,
    32'h00001888,
    32'h05000040,
    32'h00001CAD,
    32'h00001A98,
    32'h0600F000,
    32'h000018A8,
    32'hE3500000,
    32'hB3E03000,
    32'hA3A03000,
    32'hE0830000,
    32'hE0200003,
    32'hE12FFF1E,
    32'hE3700107,
    32'h82800103,
    32'h83A02205,
    32'h93A02201,
    32'h83A03801,
    32'h93A03000,
    32'hE1500002,
    32'h23833902,
    32'h20620000,
    32'hE2832A02,
    32'hE1A02682,
    32'hE1500002,
    32'h23833901,
    32'h20620000,
    32'hE2832A01,
    32'hE1A02602,
    32'hE1500002,
    32'h23833A02,
    32'h20620000,
    32'hE2832B02,
    32'hE1A02582,
    32'hE1500002,
    32'h23833A01,
    32'h20620000,
    32'hE2832B01,
    32'hE1A02502,
    32'hE1500002,
    32'h23833B02,
    32'h20620000,
    32'hE2832C02,
    32'hE1A02482,
    32'hE1500002,
    32'h23833B01,
    32'h20620000,
    32'hE2832C01,
    32'hE1A02402,
    32'hE1500002,
    32'h23833C02,
    32'h20620000,
    32'hE2832080,
    32'hE1A02382,
    32'hE1500002,
    32'h23833C01,
    32'h20620000,
    32'hE2832040,
    32'hE1A02302,
    32'hE1500002,
    32'h23833080,
    32'h20620000,
    32'hE2832020,
    32'hE1A02282,
    32'hE1500002,
    32'h23833040,
    32'h20620000,
    32'hE2832010,
    32'hE1A02202,
    32'hE1500002,
    32'h23833020,
    32'h20620000,
    32'hE2832008,
    32'hE1A02182,
    32'hE1500002,
    32'h23833010,
    32'h20620000,
    32'hE2832004,
    32'hE1A02102,
    32'hE1500002,
    32'h23833008,
    32'h20620000,
    32'hE2832002,
    32'hE1A02082,
    32'hE1500002,
    32'h23833004,
    32'h20620000,
    32'hE2832001,
    32'hE1500002,
    32'h23833002,
    32'hE1A000A3,
    32'hE12FFF1E,
    32'hE3A03301,
    32'hE5C30301,
    32'hE12FFF1E,
    32'hE3A02000,
    32'hE3A03301,
    32'hE5C32301,
    32'hE12FFF1E,
    32'hE3E0207F,
    32'hE3A03301,
    32'hE5C32301,
    32'hE12FFF1E,
    32'hE3A01000,
    32'hE3A03F82,
    32'hE3A02301,
    32'hE18210B3,
    32'hE3E0233F,
    32'hE15230B7,
    32'hE0130000,
    32'h10203003,
    32'h114230B7,
    32'hE3A01001,
    32'hE3A03F82,
    32'hE3A02301,
    32'hE20000FF,
    32'hE18210B3,
    32'hE12FFF1E,
    32'hE3500000,
    32'h01A01801,
    32'hE92D00F0,
    32'h01A00821,
    32'h0A00000E,
    32'hE3A00000,
    32'hE3A03F82,
    32'hE3A02301,
    32'hE18200B3,
    32'hE3E0233F,
    32'hE15230B7,
    32'hE1A01801,
    32'hE1A00821,
    32'hE0101003,
    32'h10213003,
    32'h114230B7,
    32'hE3A01001,
    32'hE3A03F82,
    32'hE3A02301,
    32'hE18210B3,
    32'hE3A05000,
    32'hE3A02301,
    32'hE3A0CF82,
    32'hE1A07005,
    32'hE3E0433F,
    32'hE3A06001,
    32'hE5C25301,
    32'hE18270BC,
    32'hE15430B7,
    32'hE0101003,
    32'hE0213003,
    32'h0A000005,
    32'hE31100FF,
    32'hE14430B7,
    32'hE18260BC,
    32'h0AFFFFF5,
    32'hE8BD00F0,
    32'hE12FFF1E,
    32'hE18260BC,
    32'hEAFFFFF1,
    32'hE3A00001,
    32'hE1A01000,
    32'hEAFFFFD4,
    32'hEAFFFF6A,
    32'hE0030090,
    32'hE1A03743,
    32'hE2633000,
    32'hE0832083,
    32'hE0622182,
    32'hE0832182,
    32'hE1A02742,
    32'hE2822E39,
    32'hE0020293,
    32'hE1A02742,
    32'hE2822E91,
    32'hE282200C,
    32'hE0020293,
    32'hE1A02742,
    32'hE2822EFB,
    32'hE2822006,
    32'hE0020293,
    32'hE1A02742,
    32'hE2822D5A,
    32'hE282202A,
    32'hE0020293,
    32'hE1A02742,
    32'hE2822D82,
    32'hE0223293,
    32'hE1A02742,
    32'hE2822DD9,
    32'hE2822011,
    32'hE0030392,
    32'hE1A03743,
    32'hE2833CA2,
    32'hE28330F9,
    32'hE0000093,
    32'hE1A00840,
    32'hE12FFF1E,
    32'hE92D4038,
    32'hE2515000,
    32'hE1A04000,
    32'h01A04840,
    32'h02040902,
    32'h0A000010,
    32'hE3540000,
    32'h0A000010,
    32'hE0242FC4,
    32'hE0422FC4,
    32'hE0253FC5,
    32'hE0433FC5,
    32'hE1520003,
    32'hCA000011,
    32'h0A00000D,
    32'hE1A01005,
    32'hE1A00704,
    32'hEB00047C,
    32'hEBFFFFCA,
    32'hE1A04845,
    32'hE2044902,
    32'hE2844901,
    32'hE0600004,
    32'hE8BD4038,
    32'hE12FFF1E,
    32'hE1A00845,
    32'hE2000902,
    32'hE2800901,
    32'hEAFFFFF9,
    32'hE3540000,
    32'hB3550000,
    32'hBAFFFFEE,
    32'hE1A00705,
    32'hE1A01004,
    32'hEB00046B,
    32'hEBFFFFB9,
    32'hE3540000,
    32'hA1A057A5,
    32'hA2055801,
    32'hB2800902,
    32'hA0800005,
    32'hEAFFFFEC,
    32'hE310040E,
    32'hE52D4004,
    32'h0A000018,
    32'hE1A03582,
    32'hE1A034A3,
    32'hE3C3360E,
    32'hE0833000,
    32'hE313040E,
    32'h0A000012,
    32'hE3C234FF,
    32'hE3120301,
    32'hE3C3360E,
    32'h1A000010,
    32'hE3120401,
    32'h1A00001E,
    32'hE3530000,
    32'h0A00000A,
    32'hE1A02000,
    32'hE0803083,
    32'hE0601001,
    32'hE3E044F1,
    32'hE1520004,
    32'h91D2C0B0,
    32'h859FC0A0,
    32'hE181C0B2,
    32'hE2822002,
    32'hE1520003,
    32'h1AFFFFF8,
    32'hE8BD0010,
    32'hE12FFF1E,
    32'hE3120401,
    32'hE3C11003,
    32'hE3C02003,
    32'h1A000015,
    32'hE3530000,
    32'h10621001,
    32'h13E0C4F1,
    32'h0AFFFFF5,
    32'hE152000C,
    32'h95920000,
    32'h859F0060,
    32'hE2533001,
    32'hE7810002,
    32'hE2822004,
    32'h1AFFFFF8,
    32'hEAFFFFED,
    32'hE350040F,
    32'h31D020B0,
    32'h259F203C,
    32'hE3530000,
    32'h0AFFFFE8,
    32'hE0813083,
    32'hE0C120B2,
    32'hE1510003,
    32'h1AFFFFFC,
    32'hEAFFFFE3,
    32'hE352040F,
    32'h35922000,
    32'h259F2018,
    32'hE3530000,
    32'h0AFFFFDE,
    32'hE2533001,
    32'hE4812004,
    32'h1AFFFFFC,
    32'hEAFFFFDA,
    32'h00001CAD,
    32'h1CAD1CAD,
    32'hE310040E,
    32'hE52D4004,
    32'h0A000017,
    32'hE1A03582,
    32'hE1A034A3,
    32'hE3C3360E,
    32'hE0833000,
    32'hE313040E,
    32'h0A000011,
    32'hE3C244FF,
    32'hE3120401,
    32'hE3C03003,
    32'hE3C11003,
    32'hE3C4460E,
    32'h0A00000D,
    32'hE353040F,
    32'h35932000,
    32'h259F2068,
    32'hE3540000,
    32'h0A000006,
    32'hE2813020,
    32'hE4812004,
    32'hE1510003,
    32'h1AFFFFFC,
    32'hE2444008,
    32'hE3540000,
    32'hCAFFFFF8,
    32'hE8BD0010,
    32'hE12FFF1E,
    32'hE3540000,
    32'h10631001,
    32'h13E0C4F1,
    32'h0AFFFFF9,
    32'hE2830020,
    32'hE153000C,
    32'h95932000,
    32'h859F201C,
    32'hE7812003,
    32'hE2833004,
    32'hE1530000,
    32'h1AFFFFF8,
    32'hE2444008,
    32'hE3540000,
    32'hCAFFFFF4,
    32'hEAFFFFED,
    32'hBAFFFFFB,
    32'hE59F0000,
    32'hE12FFF1E,
    32'hBAAE187F,
    32'hE3520000,
    32'hE92D0FF0,
    32'hE2422001,
    32'h0A000037,
    32'hE2800014,
    32'hE2811010,
    32'hE150C0B4,
    32'hE1A0C42C,
    32'hE28C3040,
    32'hE59F40CC,
    32'hE20330FF,
    32'hE1A03083,
    32'hE15060F8,
    32'hE19430F3,
    32'hE0040693,
    32'hE59F70B4,
    32'hE1A0C08C,
    32'hE15080F6,
    32'hE19750FC,
    32'hE00C0895,
    32'hE15070BC,
    32'hE1A04744,
    32'hE0030398,
    32'hE0050596,
    32'hE1A07807,
    32'hE1A0A804,
    32'hE1A07847,
    32'hE1A0A84A,
    32'hE00A0A97,
    32'hE1A0C74C,
    32'hE15060BA,
    32'hE1A0B80C,
    32'hE1A03743,
    32'hE1A0B84B,
    32'hE1A05745,
    32'hE00B0B97,
    32'hE1A06806,
    32'hE5107014,
    32'hE1A09803,
    32'hE1A06846,
    32'hE1A08805,
    32'hE1A09849,
    32'hE06AA007,
    32'hE0090996,
    32'hE1A08848,
    32'hE026A698,
    32'hE5107010,
    32'hE2422001,
    32'hE06B7007,
    32'hE2655000,
    32'hE0697007,
    32'hE3720001,
    32'hE14141B0,
    32'hE14150BE,
    32'hE141C0BC,
    32'hE14130BA,
    32'hE90100C0,
    32'hE2800014,
    32'hE2811010,
    32'h1AFFFFC9,
    32'hE8BD0FF0,
    32'hE12FFF1E,
    32'h00002150,
    32'hE3520000,
    32'hE92D07F0,
    32'hE2422001,
    32'h0A000021,
    32'hE1A07083,
    32'hE59FA084,
    32'hE0878083,
    32'hE2800008,
    32'hE0813003,
    32'hE150C0B4,
    32'hE1A0C42C,
    32'hE28C4040,
    32'hE20440FF,
    32'hE1A0C08C,
    32'hE15060F8,
    32'hE19A50FC,
    32'hE1A0C084,
    32'hE19AC0FC,
    32'hE15040F6,
    32'hE0090596,
    32'hE006069C,
    32'hE0050594,
    32'hE00C0C94,
    32'hE1A09749,
    32'hE2422001,
    32'hE1A06746,
    32'hE2699000,
    32'hE1A05745,
    32'hE1A0C74C,
    32'hE3720001,
    32'hE1C160B0,
    32'hE2800008,
    32'hE1C390B0,
    32'hE18150B7,
    32'hE183C0B7,
    32'hE0811008,
    32'hE0833008,
    32'h1AFFFFE2,
    32'hE8BD07F0,
    32'hE12FFF1E,
    32'h00002150,
    32'hE92D0FF0,
    32'hE310040E,
    32'hE24DD008,
    32'hE1D2C0B0,
    32'h0A000027,
    32'hE08CC000,
    32'hE31C040E,
    32'h0A000024,
    32'hE5D27002,
    32'hE3A050FF,
    32'hE2673008,
    32'hE1A05355,
    32'hE5923004,
    32'hE3A06000,
    32'hE5D2B003,
    32'hE150000C,
    32'hE1A02FA3,
    32'hE3C33102,
    32'hE58D2000,
    32'hE58D3004,
    32'hE1A0A006,
    32'h0A000016,
    32'hE4D04001,
    32'hE1A02005,
    32'hE3A03000,
    32'hE59D8000,
    32'hE0029004,
    32'hE3590000,
    32'h13888001,
    32'hE3580000,
    32'hE1A08339,
    32'h159D9004,
    32'h10888009,
    32'hE18AA618,
    32'hE086600B,
    32'hE356001F,
    32'hC3A06000,
    32'hE0833007,
    32'hC481A004,
    32'hC1A0A006,
    32'hE3530007,
    32'hE1A02712,
    32'hDAFFFFED,
    32'hE150000C,
    32'h1AFFFFE8,
    32'hE28DD008,
    32'hE8BD0FF0,
    32'hE12FFF1E,
    32'hE4902004,
    32'hE310040E,
    32'hE92D01F0,
    32'h0A00001C,
    32'hE1A02422,
    32'hE3C234FF,
    32'hE3C3360E,
    32'hE0833000,
    32'hE313040E,
    32'h0A000016,
    32'hE3520000,
    32'h0A000014,
    32'hE5D04000,
    32'hE3540000,
    32'hE280C001,
    32'h0A000012,
    32'hE3A08008,
    32'hE3140080,
    32'h1A00001A,
    32'hE5DC3000,
    32'hE2522001,
    32'hE2810001,
    32'hE28CC001,
    32'hE5C13000,
    32'h0A000007,
    32'hE1A01000,
    32'hE1A04084,
    32'hE2588001,
    32'hE20440FF,
    32'h1AFFFFF2,
    32'hE3520000,
    32'hE1A0000C,
    32'hCAFFFFEA,
    32'hE8BD01F0,
    32'hE12FFF1E,
    32'hE2804009,
    32'hE1A0000C,
    32'hE4D03001,
    32'hE2522001,
    32'hE4C13001,
    32'h0AFFFFF7,
    32'hE1500004,
    32'h1AFFFFF9,
    32'hE3520000,
    32'hCAFFFFDE,
    32'hEAFFFFF2,
    32'hE5DC0000,
    32'hE5DC3001,
    32'hE1833400,
    32'hE1A03803,
    32'hE1A07E23,
    32'hE2416001,
    32'hE1A03203,
    32'hE2420001,
    32'hE0466A23,
    32'hE2877003,
    32'hE1A05000,
    32'hE3A03000,
    32'hEA000000,
    32'hE2400001,
    32'hE7D32006,
    32'hE1530005,
    32'hE4C12001,
    32'hE2833001,
    32'hE1A02000,
    32'h0AFFFFDE,
    32'hE1570003,
    32'hCAFFFFF6,
    32'hE28CC002,
    32'hEAFFFFD3,
    32'hE92D0FF0,
    32'hE4905004,
    32'hE3520000,
    32'h01A05425,
    32'h0A000007,
    32'hE310040E,
    32'h0A000024,
    32'hE1A05425,
    32'hE3C534FF,
    32'hE3C3360E,
    32'hE0833000,
    32'hE313040E,
    32'h0A00001E,
    32'hE3550000,
    32'h0A00001C,
    32'hE3A03000,
    32'hE1A0C003,
    32'hE1A04003,
    32'hE5D07000,
    32'hE3570000,
    32'hE2806001,
    32'h0A000017,
    32'hE3A0B008,
    32'hE3170080,
    32'h1A000026,
    32'hE5D62000,
    32'hE1833C12,
    32'hE3540001,
    32'h00C130B2,
    32'h03A03000,
    32'h128CC008,
    32'h13A04001,
    32'h01A0C003,
    32'h01A04003,
    32'hE2555001,
    32'hE2866001,
    32'h0A000006,
    32'hE1A07087,
    32'hE25BB001,
    32'hE20770FF,
    32'h1AFFFFED,
    32'hE3550000,
    32'hE1A00006,
    32'hCAFFFFE5,
    32'hE8BD0FF0,
    32'hE12FFF1E,
    32'hE2807009,
    32'hE1A00006,
    32'hE4D02001,
    32'hE1833C12,
    32'hE3540001,
    32'h00C130B2,
    32'h03A03000,
    32'h128CC008,
    32'h13A04001,
    32'h01A0C003,
    32'h01A04003,
    32'hE2555001,
    32'h0AFFFFF0,
    32'hE1500007,
    32'h1AFFFFF2,
    32'hE3550000,
    32'hCAFFFFD2,
    32'hEAFFFFEB,
    32'hE5D60000,
    32'hE5D62001,
    32'hE1822400,
    32'hE1A02802,
    32'hE241A001,
    32'hE1A09E22,
    32'hE08AA004,
    32'hE1A02202,
    32'hE2450001,
    32'hE04AAA22,
    32'hE2899003,
    32'hE1A08000,
    32'hE3A02000,
    32'hEA000000,
    32'hE2400001,
    32'hE7D2500A,
    32'hE1833C15,
    32'hE3540001,
    32'h00C130B2,
    32'h03A03000,
    32'h128CC008,
    32'h13A04001,
    32'h01A0C003,
    32'h01A04003,
    32'hE1520008,
    32'hE1A05000,
    32'hE2822001,
    32'h0AFFFFCF,
    32'hE1590002,
    32'hCAFFFFEF,
    32'hE2866002,
    32'hEAFFFFC4,
    32'hE3A02001,
    32'hEAFFFF9D,
    32'hE92D0FF0,
    32'hE1A03000,
    32'hE4934004,
    32'hE24DD010,
    32'hE313040E,
    32'hE58D1000,
    32'h0A000033,
    32'hE1A02424,
    32'hE3C214FF,
    32'hE3C1160E,
    32'hE0813003,
    32'hE313040E,
    32'h0A00002D,
    32'hE5D0C004,
    32'hE2806005,
    32'hE28CC001,
    32'hE204400F,
    32'hE086C08C,
    32'hE3540008,
    32'hE51C3001,
    32'hE5D07005,
    32'hE28CC003,
    32'h0A000048,
    32'hE3520000,
    32'hDA000021,
    32'hE3A08000,
    32'hE58D800C,
    32'hE58D8004,
    32'hE58D8008,
    32'hE1A05007,
    32'hE1A09008,
    32'hE3A01102,
    32'hE3A04001,
    32'hE1110003,
    32'h11A05325,
    32'h1084B000,
    32'h1205A001,
    32'h01A0A3A5,
    32'h15DB5006,
    32'h07D45006,
    32'hE35A0000,
    32'h0A000005,
    32'hE3590000,
    32'h1A000011,
    32'hE1888005,
    32'hE3A09004,
    32'hE1A05007,
    32'hE3A04000,
    32'hE1B010A1,
    32'h049C3004,
    32'h03A01102,
    32'hE3520000,
    32'hDA000005,
    32'hE3540000,
    32'h0AFFFFE8,
    32'hE205A03F,
    32'hE28AA001,
    32'hE084408A,
    32'hEAFFFFE5,
    32'hE28DD010,
    32'hE8BD0FF0,
    32'hE12FFF1E,
    32'hE2899004,
    32'hE3590008,
    32'hE1888205,
    32'h13A04000,
    32'h11A05007,
    32'h1AFFFFEB,
    32'hE59D5004,
    32'hE2855001,
    32'hE59D400C,
    32'hE58D5004,
    32'hE3550004,
    32'hE59D5008,
    32'hE1844518,
    32'hE3A08000,
    32'hE58D400C,
    32'h0A000005,
    32'hE2855008,
    32'hE58D5008,
    32'hE1A09008,
    32'hE1A05007,
    32'hE1A04008,
    32'hEAFFFFDB,
    32'hE59D5000,
    32'hE59D400C,
    32'hE4854004,
    32'hE2422004,
    32'hE58D5000,
    32'hE1A09008,
    32'hE1A05007,
    32'hE58D800C,
    32'hE58D8004,
    32'hE58D8008,
    32'hE1A04008,
    32'hEAFFFFCF,
    32'hE3520000,
    32'hDAFFFFD8,
    32'hE3A0A000,
    32'hE1A05007,
    32'hE3A01102,
    32'hE1A0B00A,
    32'hE1A0900A,
    32'hE3A04001,
    32'hE1130001,
    32'h11A08325,
    32'h01A083A5,
    32'h10845000,
    32'h12088001,
    32'h15D55006,
    32'h07D45006,
    32'hE3580000,
    32'h0A000006,
    32'hE2899001,
    32'hE3590004,
    32'hE18AAB15,
    32'h0A00000D,
    32'hE28BB008,
    32'hE1A05007,
    32'hE3A04000,
    32'hE1B010A1,
    32'h049C3004,
    32'h03A01102,
    32'hE3520000,
    32'hDAFFFFBD,
    32'hE3540000,
    32'h0AFFFFE7,
    32'hE205803F,
    32'hE2888001,
    32'hE0844088,
    32'hEAFFFFE4,
    32'hE59D4000,
    32'hE484A004,
    32'hE3A0A000,
    32'hE58D4000,
    32'hE2422004,
    32'hE1A05007,
    32'hE1A0900A,
    32'hE1A0B00A,
    32'hE1A0400A,
    32'hEAFFFFEA,
    32'hE4902004,
    32'hE310040E,
    32'hE92D0030,
    32'h0A000017,
    32'hE1A02422,
    32'hE3C234FF,
    32'hE3C3360E,
    32'hE0833000,
    32'hE313040E,
    32'h0A000011,
    32'hE3520000,
    32'h0A00000F,
    32'hE5D04000,
    32'hE3140080,
    32'hE280C001,
    32'hE204407F,
    32'h01A03001,
    32'h1A00000B,
    32'hE4DC0001,
    32'hE4C30001,
    32'hE2522001,
    32'hE0610003,
    32'h0A000004,
    32'hE1540000,
    32'hAAFFFFF8,
    32'hE1A01003,
    32'hE1A0000C,
    32'hEAFFFFEF,
    32'hE8BD0030,
    32'hE12FFF1E,
    32'hE5D05001,
    32'hE2844003,
    32'hE1A03001,
    32'hE4C35001,
    32'hE2522001,
    32'hE061C003,
    32'h0AFFFFF6,
    32'hE154000C,
    32'hCAFFFFF9,
    32'hE280C002,
    32'hEAFFFFEF,
    32'hE92D05F0,
    32'hE2806004,
    32'hE316040E,
    32'hE3C00003,
    32'hE5900000,
    32'h0A000021,
    32'hE1A00420,
    32'hE3C034FF,
    32'hE3C3360E,
    32'hE0833006,
    32'hE313040E,
    32'h0A00001B,
    32'hE3500000,
    32'h0A000019,
    32'hE3A03000,
    32'hE1A02003,
    32'hE1A04003,
    32'hE5D67000,
    32'hE3170080,
    32'hE2865001,
    32'hE207707F,
    32'h03A0C000,
    32'h1A000012,
    32'hE4D56001,
    32'hE1833216,
    32'hE3540001,
    32'h00C130B2,
    32'h03A03000,
    32'h12822008,
    32'h13A04001,
    32'h01A02003,
    32'h01A04003,
    32'hE2500001,
    32'hE28CC001,
    32'h0A000004,
    32'hE157000C,
    32'hAAFFFFF1,
    32'hE1A06005,
    32'hE3500000,
    32'hCAFFFFE8,
    32'hE8BD05F0,
    32'hE12FFF1E,
    32'hE2405001,
    32'hE5D6A001,
    32'hE2877003,
    32'hE1A08005,
    32'hE3A0C000,
    32'hEA000000,
    32'hE2455001,
    32'hE183321A,
    32'hE3540001,
    32'h00C130B2,
    32'h03A03000,
    32'h12822008,
    32'h13A04001,
    32'h01A02003,
    32'h01A04003,
    32'hE15C0008,
    32'hE1A00005,
    32'hE28CC001,
    32'h0AFFFFEA,
    32'hE157000C,
    32'hCAFFFFF0,
    32'hE2866002,
    32'hEAFFFFE4,
    32'hE1A02000,
    32'hE492C004,
    32'hE312040E,
    32'h012FFF1E,
    32'hE1A0C42C,
    32'hE3CC34FF,
    32'hE3C3360E,
    32'hE0833002,
    32'hE313040E,
    32'h012FFF1E,
    32'hE5D03004,
    32'hE35C0001,
    32'hE2800005,
    32'hE5C13000,
    32'hD12FFF1E,
    32'hE082C00C,
    32'hE4D02001,
    32'hE0833002,
    32'hE20330FF,
    32'hE150000C,
    32'hE5E13001,
    32'h1AFFFFF9,
    32'hE12FFF1E,
    32'hE1A03000,
    32'hE92D0070,
    32'hE4936004,
    32'hE313040E,
    32'h0A00001C,
    32'hE1A06426,
    32'hE3C624FF,
    32'hE3C2260E,
    32'hE0823003,
    32'hE313040E,
    32'h0A000016,
    32'hE5D03004,
    32'hE3560001,
    32'hE2800005,
    32'hE1A0C003,
    32'hDA000011,
    32'hE3A04001,
    32'hE3A02008,
    32'hE4D05001,
    32'hE0833005,
    32'hE20330FF,
    32'hE18CC213,
    32'hE3540001,
    32'hE1A0C80C,
    32'h03A04000,
    32'hE1A0C82C,
    32'h02466002,
    32'h00C1C0B2,
    32'h12822008,
    32'h13A04001,
    32'h01A02004,
    32'h01A0C004,
    32'hE3560001,
    32'hCAFFFFEF,
    32'hE8BD0070,
    32'hE12FFF1E,
    32'hE1A03000,
    32'hE493C004,
    32'hE313040E,
    32'h012FFF1E,
    32'hE1A0C42C,
    32'hE3CC24FF,
    32'hE3C2260E,
    32'hE0823003,
    32'hE313040E,
    32'h012FFF1E,
    32'hE1D030B4,
    32'hE35C0003,
    32'hE2802006,
    32'hE1C130B0,
    32'hD12FFF1E,
    32'hE24CC004,
    32'hE2800008,
    32'hE3CCC001,
    32'hE080C00C,
    32'hE0D200B2,
    32'hE0833000,
    32'hE1A03803,
    32'hE1A03823,
    32'hE152000C,
    32'hE1E130B2,
    32'h1AFFFFF8,
    32'hE12FFF1E,
    32'hE35100B2,
    32'hE92D4038,
    32'hE59F3064,
    32'h83A010B2,
    32'hE1A05000,
    32'h92810001,
    32'hE0831001,
    32'hE5D1C200,
    32'hE20C100F,
    32'hE0831101,
    32'hE59142B4,
    32'hE1A0C22C,
    32'hE1A04C34,
    32'h83A000B3,
    32'hE0831000,
    32'hE5D1C200,
    32'hE20C100F,
    32'hE0833101,
    32'hE59302B4,
    32'h83A024FF,
    32'hE1A0C22C,
    32'hE1A01002,
    32'hE0640C30,
    32'hEBFFFBBD,
    32'hE5951004,
    32'hE0840000,
    32'hEBFFFBBA,
    32'hE8BD4038,
    32'hE12FFF1E,
    32'h00002150,
    32'hE59F325C,
    32'hE92D47F0,
    32'hE5934FF0,
    32'hE59F3254,
    32'hE5942000,
    32'hE1520003,
    32'h0A000001,
    32'hE8BD47F0,
    32'hE12FFF1E,
    32'hE5943020,
    32'hE59F223C,
    32'hE3530000,
    32'hE5842000,
    32'h15940024,
    32'h11A0E00F,
    32'h112FFF13,
    32'hE5943028,
    32'hE3530000,
    32'h15940024,
    32'h11A0E00F,
    32'h112FFF13,
    32'hE5D42004,
    32'hE3520000,
    32'hE2843E35,
    32'hE5940010,
    32'h0A000076,
    32'hE5D4100B,
    32'hE2811001,
    32'hE0621001,
    32'hE20110FF,
    32'hE0213190,
    32'hE5D46005,
    32'hE3560000,
    32'h02812E63,
    32'h01A08001,
    32'h0A000018,
    32'hE3520002,
    32'h0A000000,
    32'hE0813000,
    32'hE2807001,
    32'hE5D1C000,
    32'hE2812E63,
    32'hE1A08001,
    32'hE0877003,
    32'hE1D290D0,
    32'hE2835E63,
    32'hE1D5A0D0,
    32'hE1A0CC0C,
    32'hE0D350D1,
    32'hE089CC4C,
    32'hE08CC00A,
    32'hE08CC005,
    32'hE00C0C96,
    32'hE1A0C4CC,
    32'hE31C0080,
    32'h128CC001,
    32'hE20CC0FF,
    32'hE1530007,
    32'hE5C2C000,
    32'hE5C1C000,
    32'h1AFFFFEE,
    32'hE1B031A0,
    32'h1A00004D,
    32'hE2810E63,
    32'hE5883000,
    32'hE281C004,
    32'hE5823000,
    32'hE2802004,
    32'hE3A03000,
    32'hE58C3000,
    32'hE28C1008,
    32'hE5823000,
    32'hE1A00003,
    32'hE58C3004,
    32'hE5823004,
    32'hE2822008,
    32'hE2811010,
    32'hE2822010,
    32'hE3A03000,
    32'hE2400001,
    32'hE3700001,
    32'hE5013010,
    32'hE5023010,
    32'hE501300C,
    32'hE502300C,
    32'hE5013008,
    32'hE5023008,
    32'hE5013004,
    32'hE5023004,
    32'hE2811010,
    32'hE2822010,
    32'h1AFFFFF2,
    32'hE5D47006,
    32'hE2846090,
    32'hE1A03006,
    32'hE1A02007,
    32'hE3A08003,
    32'hE3A05000,
    32'hE5531040,
    32'hE31100C7,
    32'hE513001C,
    32'h0A00001E,
    32'hE3110080,
    32'h1A00001C,
    32'hE3110040,
    32'hE280C010,
    32'h0A000019,
    32'hE5438040,
    32'hE503C018,
    32'hE590000C,
    32'hE5030028,
    32'hE553003C,
    32'hE31100C0,
    32'h03A0C003,
    32'h13A0C013,
    32'hE35000FF,
    32'hE1A0100C,
    32'h024C1001,
    32'h020110FF,
    32'hE5435037,
    32'hE543C040,
    32'hE5035024,
    32'h05431040,
    32'hE5430037,
    32'hE5D40007,
    32'hE0211190,
    32'hE553003E,
    32'hE1A01201,
    32'hE0010190,
    32'hE1A01421,
    32'hE20110FF,
    32'hE5431036,
    32'hE5431035,
    32'hE2422001,
    32'hE20220FF,
    32'hE35200FF,
    32'hE2833040,
    32'h1AFFFFD7,
    32'hE59F3038,
    32'hE7863307,
    32'hEAFFFF79,
    32'hE1B00220,
    32'h1AFFFFBC,
    32'hE1A0C001,
    32'hEAFFFFB2,
    32'hE5D46005,
    32'hE3560000,
    32'h01A08003,
    32'h02842D26,
    32'h01A01003,
    32'h0AFFFFA5,
    32'hE1A01003,
    32'hEAFFFF8C,
    32'h03007000,
    32'h68736D53,
    32'h68736D54,
    32'hE12FFF1E,
    32'hE12FFF1E,
    32'hE59F2010,
    32'hE2803090,
    32'hE4802004,
    32'hE1500003,
    32'h1AFFFFFC,
    32'hE12FFF1E,
    32'h0000015C,
    32'hE92D4010,
    32'hE3A03000,
    32'hE24DD008,
    32'hE58D3004,
    32'hE3A02080,
    32'hE3A03301,
    32'hE2504000,
    32'hE1C320B0,
    32'h0A000064,
    32'hE3140001,
    32'h1A00006C,
    32'hE3140002,
    32'h1A000070,
    32'hE3140004,
    32'h1A000074,
    32'hE3140008,
    32'h1A000078,
    32'hE3140010,
    32'h1A00005D,
    32'hE3140080,
    32'h0A000020,
    32'hE59F31E8,
    32'hE59F11E8,
    32'hE3A02000,
    32'hE1E320B2,
    32'hE1530001,
    32'h1AFFFFFC,
    32'hE59F11D8,
    32'hE3A03381,
    32'hE3A02000,
    32'hE1E320B2,
    32'hE1530001,
    32'h1AFFFFFC,
    32'hE59F31C4,
    32'hE59F11C4,
    32'hE3A02000,
    32'hE1E320B2,
    32'hE1530001,
    32'h1AFFFFFC,
    32'hE59F31B4,
    32'hE59F11B4,
    32'hE3A02000,
    32'hE1E320B2,
    32'hE1530001,
    32'h1AFFFFFC,
    32'hE3A03301,
    32'hE3A02C01,
    32'hE3A01E13,
    32'hE3A00000,
    32'hE18300B1,
    32'hE1C322B0,
    32'hE1C323B0,
    32'hE1C322B6,
    32'hE1C323B6,
    32'hE3140020,
    32'h0A000022,
    32'hE3A03301,
    32'hE3A02000,
    32'hE3A01E11,
    32'hE18320B1,
    32'hE2811002,
    32'hE18320B1,
    32'hE3A01F45,
    32'hE18320B1,
    32'hE2811002,
    32'hE18320B1,
    32'hE3A01F46,
    32'hE18320B1,
    32'hE2811002,
    32'hE18320B1,
    32'hE3A01F47,
    32'hE18320B1,
    32'hE2811002,
    32'hE18320B1,
    32'hE3A00902,
    32'hE3A01F4D,
    32'hE18300B1,
    32'hE3A01D05,
    32'hE18320B1,
    32'hE2811002,
    32'hE18320B1,
    32'hE3A01F51,
    32'hE18320B1,
    32'hE2811002,
    32'hE18320B1,
    32'hE3A01F52,
    32'hE18320B1,
    32'hE2811002,
    32'hE18320B1,
    32'hE3A01F53,
    32'hE18320B1,
    32'hE3140040,
    32'h0A000010,
    32'hE3A03301,
    32'hE1D318B8,
    32'hE59F00DC,
    32'hE3A02000,
    32'hE3C11B3F,
    32'hE5830080,
    32'hE1C318B8,
    32'hE5C32070,
    32'hE1C329B0,
    32'hE1C329B2,
    32'hE1C329B4,
    32'hE1C329B6,
    32'hE1C329B8,
    32'hE1C329BA,
    32'hE1C329BC,
    32'hE1C329BE,
    32'hE5C32084,
    32'hE28DD008,
    32'hE8BD4010,
    32'hE12FFF1E,
    32'hE28D0004,
    32'hE3A01407,
    32'hE59F2090,
    32'hEBFFFC09,
    32'hE3140080,
    32'h0AFFFFBE,
    32'hEAFFFF9C,
    32'hE28D0004,
    32'hE3A01402,
    32'hE59F2078,
    32'hEBFFFC02,
    32'hE3140002,
    32'h0AFFFF8E,
    32'hE28D0004,
    32'hE3A01403,
    32'hE59F2064,
    32'hEBFFFBFC,
    32'hE3140004,
    32'h0AFFFF8A,
    32'hE28D0004,
    32'hE3A01405,
    32'hE59F2044,
    32'hEBFFFBF6,
    32'hE3140008,
    32'h0AFFFF86,
    32'hE28D0004,
    32'hE3A01406,
    32'hE59F2038,
    32'hEBFFFBF0,
    32'hE3140010,
    32'h0AFFFF82,
    32'hEAFFFFDF,
    32'h040001FE,
    32'h0400021E,
    32'h04000020,
    32'h0400001E,
    32'h0400005E,
    32'h040000AE,
    32'h040000DE,
    32'h880E0000,
    32'h01000100,
    32'h01010000,
    32'h01001F80,
    32'h01006000,
    32'hE1A03000,
    32'hE1A00001,
    32'hE1A01003,
    32'hEAFFFFFF,
    32'hE210C102,
    32'h42600000,
    32'hE2113102,
    32'h42611000,
    32'hE02CC003,
    32'hE3A02000,
    32'hE3A03001,
    32'hE1510000,
    32'h91A01081,
    32'h91A03083,
    32'h9AFFFFFB,
    32'hE1500001,
    32'h20400001,
    32'h21822003,
    32'hE1B030A3,
    32'h31A010A1,
    32'h3AFFFFF9,
    32'hE1A01000,
    32'hE1A03002,
    32'hE1A00002,
    32'hE31C0102,
    32'h42600000,
    32'hE12FFF1E,
    32'hE3A03301,
    32'hE5532006,
    32'hEB000007,
    32'hE3520000,
    32'hE9131FFF,
    32'h13A0E402,
    32'h03A0E302,
    32'hE3A0001F,
    32'hE129F000,
    32'hE3A00000,
    32'hE12FFF1E,
    32'hE3A000D3,
    32'hE129F000,
    32'hE59FD044,
    32'hE3A0E000,
    32'hE169F00E,
    32'hE3A000D2,
    32'hE129F000,
    32'hE59FD02C,
    32'hE3A0E000,
    32'hE169F00E,
    32'hE3A0005F,
    32'hE129F000,
    32'hE59FD014,
    32'hE3B00000,
    32'hE2501C02,
    32'hE7830001,
    32'hE2911004,
    32'hBAFFFFFC,
    32'hE12FFF1E,
    32'h03007F00,
    32'h03007FA0,
    32'h03007FE0,
    32'h04210000,
    32'h0C630842,
    32'h18C61084,
    32'h21081CE7,
    32'h2D6B294A,
    32'h63184631,
    32'h77BD6F7B,
    32'h7FFF7BDE,
    32'h00080010,
    32'hF000003F,
    32'hF001F001,
    32'hF001F001,
    32'hFF01F001,
    32'h01F001F0,
    32'h01F001F0,
    32'h01F001F0,
    32'h01F001F0,
    32'hF001F0FF,
    32'hF001F001,
    32'hF001F001,
    32'h7001F001,
    32'h00011D07,
    32'hF001F002,
    32'h030B4001,
    32'h040140A0,
    32'h06000500,
    32'h01F00700,
    32'h4001F0C1,
    32'h0900080B,
    32'h84400A00,
    32'h0C000B00,
    32'h0E000D00,
    32'h000F0600,
    32'hF0110010,
    32'h1205A098,
    32'h00130002,
    32'h00150014,
    32'h00081619,
    32'h20180017,
    32'h1A001921,
    32'h1B290080,
    32'h1D001C00,
    32'h00001E00,
    32'h0020001F,
    32'h00220021,
    32'h24002300,
    32'h26002500,
    32'h00270000,
    32'h00290028,
    32'h2B00002A,
    32'h2D002C00,
    32'h00002E00,
    32'h0030002F,
    32'h88320031,
    32'h00335B00,
    32'h35612034,
    32'h20803600,
    32'h3800373F,
    32'h3A003900,
    32'h003B0000,
    32'h003D003C,
    32'h3F00003E,
    32'h41004000,
    32'h00004200,
    32'h00440043,
    32'h00460045,
    32'h48004700,
    32'h4A004900,
    32'h004B0008,
    32'h4D99204C,
    32'h20804E00,
    32'h50004FA1,
    32'h52005100,
    32'h00530000,
    32'h00550054,
    32'h57000056,
    32'h59005800,
    32'h00005A00,
    32'h005C005B,
    32'h005E005D,
    32'h60005F00,
    32'h62006100,
    32'h00630000,
    32'h00650064,
    32'h67000866,
    32'hD9006800,
    32'h206A0069,
    32'hE1406B00,
    32'h006D006C,
    32'h6F00386E,
    32'h01F001F0,
    32'h00700B40,
    32'h72002071,
    32'h00731F81,
    32'hE3750074,
    32'h01F001F0,
    32'h00760B40,
    32'hF05DF177,
    32'h01F0FF01,
    32'h01F001F0,
    32'h01F001F0,
    32'h01F001F0,
    32'hF0FF01F0,
    32'hF001F001,
    32'hF001F001,
    32'hF001F001,
    32'hFF01F001,
    32'h01F001F0,
    32'h01F001F0,
    32'h01F001F0,
    32'h01F001F0,
    32'hF001F0FF,
    32'hF001F001,
    32'hF001F001,
    32'hF001F001,
    32'h01F0FF01,
    32'h01F001F0,
    32'h01F001F0,
    32'h01F001F0,
    32'hF0FF01F0,
    32'hF001F001,
    32'hF001F001,
    32'hF001F001,
    32'hFF01F001,
    32'h01F001F0,
    32'h01F001F0,
    32'h01F001F0,
    32'h01F001F0,
    32'hF001F0FE,
    32'hF001F001,
    32'hF001F001,
    32'h00016001,
    32'h000F0010,
    32'hF000003C,
    32'hF001F001,
    32'h410D1001,
    32'h88883376,
    32'h077015F0,
    32'h1FF08888,
    32'h78101FA0,
    32'h15F00247,
    32'h00009200,
    32'h00DA2000,
    32'h00FFA300,
    32'hFFEA2020,
    32'h00951F00,
    32'h00EDB940,
    32'hFFFEB910,
    32'hFFFFFEB7,
    32'hFFFFFD14,
    32'h00EF0110,
    32'h06FFAB06,
    32'hBA14ADFF,
    32'h901030ED,
    32'hAB0CCD05,
    32'h40275699,
    32'hFF1DF058,
    32'h555508FF,
    32'h77505555,
    32'hC0BDEFFF,
    32'h23B04700,
    32'hEDCA9995,
    32'h10280000,
    32'h179B10A5,
    32'h5ACEA000,
    32'hFF000901,
    32'h4B004ACF,
    32'h7E0029CE,
    32'h7F10AE56,
    32'h938700EB,
    32'hBFD00400,
    32'hD000A703,
    32'hCFD4005B,
    32'h107B0005,
    32'hA801F008,
    32'h00300E10,
    32'h17007013,
    32'h85A200B0,
    32'hFFD94300,
    32'hD80060FF,
    32'h80DB00B1,
    32'hFBAE0A00,
    32'hFE3BFFFF,
    32'h04DF00FF,
    32'h00AFFFFF,
    32'h0401BDFF,
    32'h003AFF00,
    32'h44008D00,
    32'h48F01862,
    32'h000001F0,
    32'hF01200D0,
    32'hA00380C2,
    32'hCDDDDD21,
    32'h1A420105,
    32'h8E4601AE,
    32'hF0BF4A01,
    32'hD0CBB03E,
    32'hDD01DB02,
    32'hFFFC0BDD,
    32'h03500CFF,
    32'h5022F0D6,
    32'h63015009,
    32'h501FE1F0,
    32'h45755509,
    32'h7DF09B01,
    32'h01400680,
    32'h3FF0A0A3,
    32'h013F60C0,
    32'h0004DF93,
    32'h09FDA200,
    32'hD91000FF,
    32'hFB402702,
    32'hC6622500,
    32'h30605741,
    32'h0203BFFF,
    32'h02A41A03,
    32'h0B029E07,
    32'h3F0204CF,
    32'hFF0BEA1A,
    32'h01B36CFF,
    32'h1000705C,
    32'h30AA59F0,
    32'hFF70010B,
    32'hE91D00D4,
    32'hC8FA0F02,
    32'h6300B601,
    32'hDB00FC40,
    32'h540000FE,
    32'h609B0260,
    32'h305C8D02,
    32'hB107DF5F,
    32'h20028F00,
    32'h00B601D3,
    32'h03309FFF,
    32'hE08BC1F5,
    32'h02CB4203,
    32'hDA02DFD5,
    32'h2A9A00BF,
    32'h9601C4BF,
    32'h209A0190,
    32'hAB1A9E11,
    32'h007D9A00,
    32'h2903BF9E,
    32'h000C00EF,
    32'hFE00006E,
    32'hFB0001BF,
    32'h003C09EF,
    32'h917B00D7,
    32'h9103F08B,
    32'h0021109F,
    32'hDBA74000,
    32'hFFFDB700,
    32'hFFFD9008,
    32'h1B64009E,
    32'hFF20FFFA,
    32'h22F95009,
    32'hFE000122,
    32'h15ABDE10,
    32'h129C5E03,
    32'hEF4CFFD9,
    32'h00FF7A01,
    32'h3E702001,
    32'h00352222,
    32'h00EF02B0,
    32'h07002A03,
    32'h600B008D,
    32'h500F10BF,
    32'h4410013F,
    32'hB80A1BFF,
    32'h039CFFFE,
    32'hA403CDA1,
    32'hFB9902BE,
    32'hA2002CFF,
    32'h00135951,
    32'hBF210000,
    32'hFFFA003A,
    32'h0003AF2D,
    32'h7A000A76,
    32'h011D7E10,
    32'h7F608553,
    32'h3AFFFF51,
    32'h11AA9A01,
    32'h03BB580B,
    32'h69003466,
    32'h00009C40,
    32'h8ABB15BA,
    32'h3AFA0301,
    32'h01EC7F13,
    32'h04B758C8,
    32'h0B044007,
    32'h4453B931,
    32'hCB920B00,
    32'h380350BC,
    32'h031F04B5,
    32'hBFFF003F,
    32'h4BFFDA99,
    32'hFD408000,
    32'h004BD951,
    32'h08DF2220,
    32'hF500D06A,
    32'h009F0300,
    32'h0B00AF07,
    32'h70D040BF,
    32'hA81002BF,
    32'hC0B66FFF,
    32'h3D011B00,
    32'hFFDBBDFF,
    32'h844837DF,
    32'h2000BF41,
    32'hABBB0C02,
    32'h4B049505,
    32'hA701119D,
    32'hCB820497,
    32'h01A08714,
    32'hAA32AE3F,
    32'hBA400345,
    32'hC8AB30CC,
    32'h9F449B04,
    32'hFEA99AFF,
    32'h1002FF0D,
    32'h141F64FA,
    32'h66024B17,
    32'hA31A0280,
    32'hFB4005CF,
    32'h019007DF,
    32'h74D80960,
    32'h0112213F,
    32'hCEEC10A6,
    32'hFF7D10AB,
    32'h709229EF,
    32'h50E301FF,
    32'h989D527F,
    32'hB3599999,
    32'h10AFFF04,
    32'hAFBB0103,
    32'h232014D7,
    32'hFFF00163,
    32'hFFFBBBB2,
    32'hF91B05F3,
    32'h13500310,
    32'h8F125E22,
    32'hBBDF9312,
    32'hFF3C5301,
    32'h500320DF,
    32'h137F2313,
    32'h0FFFA063,
    32'hFFDBBBA0,
    32'h0320DE01,
    32'h7F131350,
    32'h206313DF,
    32'h3F20EF03,
    32'h1340AA42,
    32'h3A437F13,
    32'h00EE049C,
    32'hA3034007,
    32'h00CC044D,
    32'h2705ACE9,
    32'hA12B05B4,
    32'h57222F05,
    32'h002AFFFE,
    32'h08033040,
    32'h030A7A03,
    32'h03AB2B7E,
    32'h86036D82,
    32'h9E8A039D,
    32'h03202731,
    32'h336753DD,
    32'hCF01506F,
    32'h87137F13,
    32'h7F3B1200,
    32'h236753E9,
    32'h2077136F,
    32'h03F303EB,
    32'h68F7331F,
    32'h8003F0BF,
    32'h6305A107,
    32'h44EFFC30,
    32'h4B830508,
    32'hCF01B200,
    32'hDF69FD50,
    32'h77065A00,
    32'h707B06B3,
    32'h564B03FF,
    32'h7C4F034C,
    32'h109C5303,
    32'h9C7F0603,
    32'h7C8206A8,
    32'h064C8606,
    32'hFFFC1C8A,
    32'hFD08EF17,
    32'h00FE0300,
    32'h20960607,
    32'h0F10EF07,
    32'hC7051710,
    32'h04E73009,
    32'h0103E0A3,
    32'h3E04A503,
    32'hEF7202EF,
    32'hBAD406B9,
    32'h10B00370,
    32'hA004EF0F,
    32'h0BFF5F13,
    32'h00B15000,
    32'h03F00003,
    32'h99990B30,
    32'hFD431319,
    32'h0B4003F0,
    32'h03076B03,
    32'h0B5003F0,
    32'hDF431310,
    32'h0B6003F0,
    32'h05F30408,
    32'h4003F065,
    32'hDD43130B,
    32'h078003F0,
    32'hF083076F,
    32'hF90B6003,
    32'hF8715F01,
    32'h03F0E500,
    32'h00000B30,
    32'h590308F5,
    32'hF10708F2,
    32'h0F0003F0,
    32'hC50419FF,
    32'hF104496A,
    32'h08691913,
    32'h2408691C,
    32'h2508B749,
    32'h027D1129,
    32'h03087F78,
    32'h0B3003F0,
    32'hD6A305BF,
    32'h03F06407,
    32'h4B930770,
    32'h5F8303F0,
    32'hA303F0FF,
    32'hC303F05F,
    32'h3603F05F,
    32'h062743DF,
    32'h00FF1C72,
    32'h15370380,
    32'h00280897,
    32'h5733FAC5,
    32'h2F132753,
    32'h27183713,
    32'h1BCE065D,
    32'h065743DA,
    32'hE413C4D9,
    32'hD6206F48,
    32'hFF25FFE9,
    32'hAF23096D,
    32'h076F0800,
    32'h04A47718,
    32'hA603AE53,
    32'h440640FF,
    32'hF8D9D800,
    32'h191717DF,
    32'h2007A713,
    32'hDFF64AFF,
    32'hB0B817E3,
    32'h4473B35F,
    32'h6CD73444,
    32'h17B60316,
    32'h9FF090B7,
    32'h100CBF29,
    32'h0CFA0903,
    32'h0C170986,
    32'hA8444443,
    32'h1B030596,
    32'hFFFEA100,
    32'hFEC9209E,
    32'h60000BEF,
    32'h6606DCBA,
    32'h04CDA733,
    32'hCF068073,
    32'hDFFEDDDF,
    32'h0DBDFF4A,
    32'h2344017A,
    32'hEF77D917,
    32'h63D3064C,
    32'h26D74607,
    32'h444430DF,
    32'h73C33FA8,
    32'h607DB0EC,
    32'h427B93BF,
    32'h73B35FB1,
    32'hCADD4444,
    32'h4473D3F2,
    32'h73D37FB0,
    32'hB843A908,
    32'h73B38CDF,
    32'hB0303444,
    32'h4473C3BF,
    32'hEBB8DA14,
    32'hC14173D3,
    32'h4073F35F,
    32'h80091FB1,
    32'h90094909,
    32'h1009FFFE,
    32'h4D089CC9,
    32'h5EB14460,
    32'h3B0BE309,
    32'h710429EF,
    32'hEDDEFFFF,
    32'h21BDAB0B,
    32'hA1444335,
    32'hAFFF039F,
    32'h0BAFAF08,
    32'h0AAF41D6,
    32'h4442AFF7,
    32'h8DB92444,
    32'hC073D3FB,
    32'hF273C37F,
    32'h2073D35E,
    32'h73C3DFB1,
    32'hC0D04470,
    32'hA71201F0,
    32'h710000C7,
    32'h2000FC03,
    32'h0B10FFD9,
    32'hAA471AAC,
    32'h0AAEDE06,
    32'hA20C5C57,
    32'h03670A0A,
    32'h2A2B08FD,
    32'hF2131777,
    32'h079F9232,
    32'hE71C100B,
    32'hEB1CA264,
    32'h8100F70C,
    32'h16BEBFAA,
    32'hADC30C96,
    32'hACF60C16,
    32'hFF1CFA1C,
    32'h040DC6A4,
    32'h20000F1D,
    32'h30EF02A7,
    32'h00872852,
    32'hAAABEF59,
    32'hDDEDDC89,
    32'h8C1FF08F,
    32'hA8A61F6A,
    32'hADD51CAA,
    32'hBA00EF2F,
    32'h0AA46C00,
    32'h1D194050,
    32'hDC09AD77,
    32'hBFFF0307,
    32'h39BD0039,
    32'hF30AC31B,
    32'hBFD808B4,
    32'hA60C8A0B,
    32'h00D0FD00,
    32'h12F0D394,
    32'h09BA0770,
    32'h7D4431CC,
    32'hC0FFF38F,
    32'h1FE0AFBD,
    32'h559ABDEF,
    32'hF1D83445,
    32'h160A40B4,
    32'h01A012F0,
    32'h01920000,
    32'h04B50323,
    32'h07D50645,
    32'h0AF10964,
    32'h0E050C7C,
    32'h11110F8C,
    32'h14131294,
    32'h1708158F,
    32'h19EF187D,
    32'h1CC61B5D,
    32'h1F8B1E2B,
    32'h223D20E7,
    32'h24DA238E,
    32'h275F261F,
    32'h29CD2899,
    32'h2C212AFA,
    32'h2E5A2D41,
    32'h30762F6B,
    32'h32743179,
    32'h34533367,
    32'h36123536,
    32'h37AF36E5,
    32'h392A3871,
    32'h3A8239DA,
    32'h3BB63B20,
    32'h3CC53C42,
    32'h3DAE3D3E,
    32'h3E713E14,
    32'h3F0E3EC5,
    32'h3F843F4E,
    32'h3FD33FB1,
    32'h3FFB3FEC,
    32'h3FFB4000,
    32'h3FD33FEC,
    32'h3F843FB1,
    32'h3F0E3F4E,
    32'h3E713EC5,
    32'h3DAE3E14,
    32'h3CC53D3E,
    32'h3BB63C42,
    32'h3A823B20,
    32'h392A39DA,
    32'h37AF3871,
    32'h361236E5,
    32'h34533536,
    32'h32743367,
    32'h30763179,
    32'h2E5A2F6B,
    32'h2C212D41,
    32'h29CD2AFA,
    32'h275F2899,
    32'h24DA261F,
    32'h223D238E,
    32'h1F8B20E7,
    32'h1CC61E2B,
    32'h19EF1B5D,
    32'h1708187D,
    32'h1413158F,
    32'h11111294,
    32'h0E050F8C,
    32'h0AF10C7C,
    32'h07D50964,
    32'h04B50645,
    32'h01920323,
    32'hFE6E0000,
    32'hFB4BFCDD,
    32'hF82BF9BB,
    32'hF50FF69C,
    32'hF1FBF384,
    32'hEEEFF074,
    32'hEBEDED6C,
    32'hE8F8EA71,
    32'hE611E783,
    32'hE33AE4A3,
    32'hE075E1D5,
    32'hDDC3DF19,
    32'hDB26DC72,
    32'hD8A1D9E1,
    32'hD633D767,
    32'hD3DFD506,
    32'hD1A6D2BF,
    32'hCF8AD095,
    32'hCD8CCE87,
    32'hCBADCC99,
    32'hC9EECACA,
    32'hC851C91B,
    32'hC6D6C78F,
    32'hC57EC626,
    32'hC44AC4E0,
    32'hC33BC3BE,
    32'hC252C2C2,
    32'hC18FC1EC,
    32'hC0F2C13B,
    32'hC07CC0B2,
    32'hC02DC04F,
    32'hC005C014,
    32'hC005C000,
    32'hC02DC014,
    32'hC07CC04F,
    32'hC0F2C0B2,
    32'hC18FC13B,
    32'hC252C1EC,
    32'hC33BC2C2,
    32'hC44AC3BE,
    32'hC57EC4E0,
    32'hC6D6C626,
    32'hC851C78F,
    32'hC9EEC91B,
    32'hCBADCACA,
    32'hCD8CCC99,
    32'hCF8ACE87,
    32'hD1A6D095,
    32'hD3DFD2BF,
    32'hD633D506,
    32'hD8A1D767,
    32'hDB26D9E1,
    32'hDDC3DC72,
    32'hE075DF19,
    32'hE33AE1D5,
    32'hE611E4A3,
    32'hE8F8E783,
    32'hEBEDEA71,
    32'hEEEFED6C,
    32'hF1FBF074,
    32'hF50FF384,
    32'hF82BF69C,
    32'hFB4BF9BB,
    32'hFE6EFCDD,
    32'hE3E2E1E0,
    32'hE7E6E5E4,
    32'hEBEAE9E8,
    32'hD3D2D1D0,
    32'hD7D6D5D4,
    32'hDBDAD9D8,
    32'hC3C2C1C0,
    32'hC7C6C5C4,
    32'hCBCAC9C8,
    32'hB3B2B1B0,
    32'hB7B6B5B4,
    32'hBBBAB9B8,
    32'hA3A2A1A0,
    32'hA7A6A5A4,
    32'hABAAA9A8,
    32'h93929190,
    32'h97969594,
    32'h9B9A9998,
    32'h83828180,
    32'h87868584,
    32'h8B8A8988,
    32'h73727170,
    32'h77767574,
    32'h7B7A7978,
    32'h63626160,
    32'h67666564,
    32'h6B6A6968,
    32'h53525150,
    32'h57565554,
    32'h5B5A5958,
    32'h43424140,
    32'h47464544,
    32'h4B4A4948,
    32'h33323130,
    32'h37363534,
    32'h3B3A3938,
    32'h23222120,
    32'h27262524,
    32'h2B2A2928,
    32'h13121110,
    32'h17161514,
    32'h1B1A1918,
    32'h03020100,
    32'h07060504,
    32'h0B0A0908,
    32'h80000000,
    32'h879C7C97,
    32'h8FACD61E,
    32'h9837F052,
    32'hA14517CC,
    32'hAADC0848,
    32'hB504F334,
    32'hBFC886BB,
    32'hCB2FF52A,
    32'hD744FCCB,
    32'hE411F03A,
    32'hF1A1BF39,
    32'h52416B64,
    32'h0000004D,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000
};

`endif